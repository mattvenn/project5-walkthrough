VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rgb_mixer
  CLASS BLOCK ;
  FOREIGN rgb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 159.840 100.000 160.440 ;
    END
  END clk
  PIN enc0_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END enc0_a
  PIN enc0_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 204.040 100.000 204.640 ;
    END
  END enc0_b
  PIN enc1_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 71.440 100.000 72.040 ;
    END
  END enc1_a
  PIN enc1_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 246.000 13.250 250.000 ;
    END
  END enc1_b
  PIN enc2_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END enc2_a
  PIN enc2_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 27.240 100.000 27.840 ;
    END
  END enc2_b
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 246.000 55.110 250.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_oeb[3]
  PIN pwm0_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 246.000 96.970 250.000 ;
    END
  END pwm0_out
  PIN pwm1_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END pwm1_out
  PIN pwm2_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END pwm2_out
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END reset
  PIN sync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 115.640 100.000 116.240 ;
    END
  END sync
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.550 10.640 21.150 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.855 10.640 80.455 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 236.725 ;
      LAYER met1 ;
        RECT 0.070 10.640 96.990 236.880 ;
      LAYER met2 ;
        RECT 0.100 245.720 12.690 246.570 ;
        RECT 13.530 245.720 54.550 246.570 ;
        RECT 55.390 245.720 96.410 246.570 ;
        RECT 0.100 4.280 96.960 245.720 ;
        RECT 0.650 4.000 41.670 4.280 ;
        RECT 42.510 4.000 83.530 4.280 ;
        RECT 84.370 4.000 96.960 4.280 ;
      LAYER met3 ;
        RECT 4.000 222.040 96.000 236.805 ;
        RECT 4.400 220.640 96.000 222.040 ;
        RECT 4.000 205.040 96.000 220.640 ;
        RECT 4.000 203.640 95.600 205.040 ;
        RECT 4.000 177.840 96.000 203.640 ;
        RECT 4.400 176.440 96.000 177.840 ;
        RECT 4.000 160.840 96.000 176.440 ;
        RECT 4.000 159.440 95.600 160.840 ;
        RECT 4.000 133.640 96.000 159.440 ;
        RECT 4.400 132.240 96.000 133.640 ;
        RECT 4.000 116.640 96.000 132.240 ;
        RECT 4.000 115.240 95.600 116.640 ;
        RECT 4.000 89.440 96.000 115.240 ;
        RECT 4.400 88.040 96.000 89.440 ;
        RECT 4.000 72.440 96.000 88.040 ;
        RECT 4.000 71.040 95.600 72.440 ;
        RECT 4.000 45.240 96.000 71.040 ;
        RECT 4.400 43.840 96.000 45.240 ;
        RECT 4.000 28.240 96.000 43.840 ;
        RECT 4.000 26.840 95.600 28.240 ;
        RECT 4.000 10.715 96.000 26.840 ;
      LAYER met4 ;
        RECT 21.550 10.640 33.970 236.880 ;
        RECT 36.370 10.640 48.800 236.880 ;
        RECT 51.200 10.640 63.625 236.880 ;
        RECT 66.025 10.640 78.455 236.880 ;
  END
END rgb_mixer
END LIBRARY

