magic
tech sky130A
magscale 1 2
timestamp 1647353466
<< viali >>
rect 11529 47209 11563 47243
rect 18061 47209 18095 47243
rect 2789 47005 2823 47039
rect 17877 47005 17911 47039
rect 2973 46937 3007 46971
rect 8953 45917 8987 45951
rect 9137 45917 9171 45951
rect 9045 45781 9079 45815
rect 6745 45509 6779 45543
rect 8125 45509 8159 45543
rect 8325 45509 8359 45543
rect 9965 45509 9999 45543
rect 7021 45441 7055 45475
rect 7481 45441 7515 45475
rect 7665 45441 7699 45475
rect 9137 45441 9171 45475
rect 9321 45441 9355 45475
rect 9873 45441 9907 45475
rect 10149 45441 10183 45475
rect 11529 45441 11563 45475
rect 11713 45441 11747 45475
rect 6745 45373 6779 45407
rect 9413 45373 9447 45407
rect 8493 45305 8527 45339
rect 10149 45305 10183 45339
rect 6929 45237 6963 45271
rect 7481 45237 7515 45271
rect 8309 45237 8343 45271
rect 8953 45237 8987 45271
rect 11529 45237 11563 45271
rect 7389 45033 7423 45067
rect 11529 44965 11563 44999
rect 5549 44829 5583 44863
rect 7573 44829 7607 44863
rect 7665 44829 7699 44863
rect 8217 44829 8251 44863
rect 8401 44829 8435 44863
rect 8953 44829 8987 44863
rect 9209 44829 9243 44863
rect 10885 44829 10919 44863
rect 11161 44829 11195 44863
rect 11437 44829 11471 44863
rect 11621 44829 11655 44863
rect 12081 44829 12115 44863
rect 5816 44761 5850 44795
rect 12173 44761 12207 44795
rect 6929 44693 6963 44727
rect 8309 44693 8343 44727
rect 10333 44693 10367 44727
rect 5733 44489 5767 44523
rect 6377 44489 6411 44523
rect 11529 44489 11563 44523
rect 7490 44421 7524 44455
rect 1869 44353 1903 44387
rect 5641 44353 5675 44387
rect 5825 44353 5859 44387
rect 8401 44353 8435 44387
rect 8677 44353 8711 44387
rect 10710 44353 10744 44387
rect 10977 44353 11011 44387
rect 12653 44353 12687 44387
rect 12909 44353 12943 44387
rect 2145 44285 2179 44319
rect 7757 44285 7791 44319
rect 8585 44217 8619 44251
rect 8217 44149 8251 44183
rect 9597 44149 9631 44183
rect 6285 43945 6319 43979
rect 8309 43945 8343 43979
rect 10333 43945 10367 43979
rect 11529 43945 11563 43979
rect 13369 43945 13403 43979
rect 6377 43877 6411 43911
rect 13277 43877 13311 43911
rect 6193 43809 6227 43843
rect 6929 43809 6963 43843
rect 11161 43809 11195 43843
rect 12265 43809 12299 43843
rect 13369 43809 13403 43843
rect 6469 43741 6503 43775
rect 7196 43741 7230 43775
rect 8953 43741 8987 43775
rect 9220 43741 9254 43775
rect 10793 43741 10827 43775
rect 10977 43741 11011 43775
rect 11069 43741 11103 43775
rect 11345 43741 11379 43775
rect 12357 43741 12391 43775
rect 13001 43673 13035 43707
rect 11989 43605 12023 43639
rect 13093 43605 13127 43639
rect 7221 43401 7255 43435
rect 9873 43401 9907 43435
rect 12449 43401 12483 43435
rect 7021 43333 7055 43367
rect 9505 43333 9539 43367
rect 9597 43333 9631 43367
rect 10333 43333 10367 43367
rect 8125 43265 8159 43299
rect 8309 43265 8343 43299
rect 9229 43265 9263 43299
rect 9377 43265 9411 43299
rect 9694 43265 9728 43299
rect 10701 43265 10735 43299
rect 10793 43265 10827 43299
rect 12081 43265 12115 43299
rect 10425 43197 10459 43231
rect 11989 43197 12023 43231
rect 7389 43129 7423 43163
rect 7205 43061 7239 43095
rect 7941 43061 7975 43095
rect 10517 43061 10551 43095
rect 9137 42857 9171 42891
rect 8953 42721 8987 42755
rect 10977 42721 11011 42755
rect 9229 42653 9263 42687
rect 9873 42653 9907 42687
rect 11069 42653 11103 42687
rect 8953 42517 8987 42551
rect 9781 42517 9815 42551
rect 9137 42313 9171 42347
rect 10333 42313 10367 42347
rect 7573 42177 7607 42211
rect 8401 42177 8435 42211
rect 8585 42177 8619 42211
rect 8769 42177 8803 42211
rect 8953 42177 8987 42211
rect 10241 42177 10275 42211
rect 10425 42177 10459 42211
rect 8677 42109 8711 42143
rect 7849 41973 7883 42007
rect 8677 41225 8711 41259
rect 8309 41157 8343 41191
rect 8125 41089 8159 41123
rect 8401 41089 8435 41123
rect 8493 41089 8527 41123
rect 14657 41089 14691 41123
rect 14841 41089 14875 41123
rect 15301 41089 15335 41123
rect 15945 41089 15979 41123
rect 18153 41089 18187 41123
rect 14473 41021 14507 41055
rect 15485 40885 15519 40919
rect 16129 40885 16163 40919
rect 17969 40885 18003 40919
rect 6837 40681 6871 40715
rect 8309 40681 8343 40715
rect 9137 40681 9171 40715
rect 7941 40477 7975 40511
rect 9229 40477 9263 40511
rect 12725 40477 12759 40511
rect 15577 40477 15611 40511
rect 16037 40477 16071 40511
rect 16293 40477 16327 40511
rect 6791 40443 6825 40477
rect 7021 40409 7055 40443
rect 8125 40409 8159 40443
rect 15332 40409 15366 40443
rect 6653 40341 6687 40375
rect 12909 40341 12943 40375
rect 14197 40341 14231 40375
rect 17417 40341 17451 40375
rect 7573 40137 7607 40171
rect 7849 40069 7883 40103
rect 12878 40069 12912 40103
rect 5641 40001 5675 40035
rect 5837 40001 5871 40035
rect 6561 40001 6595 40035
rect 7732 40001 7766 40035
rect 7941 40001 7975 40035
rect 8124 40001 8158 40035
rect 8217 40001 8251 40035
rect 10517 40001 10551 40035
rect 11989 40001 12023 40035
rect 12173 40001 12207 40035
rect 15016 40001 15050 40035
rect 16865 40001 16899 40035
rect 6837 39933 6871 39967
rect 10425 39933 10459 39967
rect 12633 39933 12667 39967
rect 14749 39933 14783 39967
rect 16681 39933 16715 39967
rect 17049 39933 17083 39967
rect 16129 39865 16163 39899
rect 5825 39797 5859 39831
rect 6377 39797 6411 39831
rect 6745 39797 6779 39831
rect 10793 39797 10827 39831
rect 12081 39797 12115 39831
rect 14013 39797 14047 39831
rect 10793 39593 10827 39627
rect 11897 39593 11931 39627
rect 12817 39593 12851 39627
rect 14749 39593 14783 39627
rect 6377 39525 6411 39559
rect 8401 39525 8435 39559
rect 10241 39525 10275 39559
rect 6837 39457 6871 39491
rect 9965 39457 9999 39491
rect 10977 39457 11011 39491
rect 11989 39457 12023 39491
rect 14565 39457 14599 39491
rect 4997 39389 5031 39423
rect 7113 39389 7147 39423
rect 8125 39389 8159 39423
rect 9873 39389 9907 39423
rect 10701 39389 10735 39423
rect 11713 39389 11747 39423
rect 11805 39389 11839 39423
rect 12449 39389 12483 39423
rect 12633 39389 12667 39423
rect 13553 39389 13587 39423
rect 14749 39389 14783 39423
rect 15577 39389 15611 39423
rect 15669 39389 15703 39423
rect 16405 39389 16439 39423
rect 16497 39389 16531 39423
rect 5264 39321 5298 39355
rect 8401 39321 8435 39355
rect 14473 39321 14507 39355
rect 15393 39321 15427 39355
rect 8217 39253 8251 39287
rect 10977 39253 11011 39287
rect 13369 39253 13403 39287
rect 14933 39253 14967 39287
rect 16221 39253 16255 39287
rect 5647 39049 5681 39083
rect 7757 39049 7791 39083
rect 8953 39049 8987 39083
rect 12081 39049 12115 39083
rect 15117 39049 15151 39083
rect 15761 39049 15795 39083
rect 9873 38981 9907 39015
rect 11897 38981 11931 39015
rect 15301 38981 15335 39015
rect 3617 38913 3651 38947
rect 3873 38913 3907 38947
rect 5549 38913 5583 38947
rect 5733 38913 5767 38947
rect 5825 38913 5859 38947
rect 6644 38913 6678 38947
rect 8217 38913 8251 38947
rect 8401 38913 8435 38947
rect 8585 38913 8619 38947
rect 8769 38913 8803 38947
rect 9597 38913 9631 38947
rect 9689 38913 9723 38947
rect 10425 38913 10459 38947
rect 10701 38913 10735 38947
rect 11713 38913 11747 38947
rect 12909 38913 12943 38947
rect 13176 38913 13210 38947
rect 14933 38913 14967 38947
rect 15025 38913 15059 38947
rect 15945 38913 15979 38947
rect 6377 38845 6411 38879
rect 8493 38845 8527 38879
rect 10517 38845 10551 38879
rect 10885 38845 10919 38879
rect 9873 38777 9907 38811
rect 10609 38777 10643 38811
rect 4997 38709 5031 38743
rect 14289 38709 14323 38743
rect 14749 38709 14783 38743
rect 12541 38505 12575 38539
rect 15485 38505 15519 38539
rect 6653 38437 6687 38471
rect 10977 38437 11011 38471
rect 7113 38369 7147 38403
rect 7389 38369 7423 38403
rect 9781 38369 9815 38403
rect 11713 38369 11747 38403
rect 14105 38369 14139 38403
rect 3801 38301 3835 38335
rect 3985 38301 4019 38335
rect 5273 38301 5307 38335
rect 9689 38301 9723 38335
rect 10793 38301 10827 38335
rect 11621 38301 11655 38335
rect 12449 38301 12483 38335
rect 12633 38301 12667 38335
rect 13369 38301 13403 38335
rect 5540 38233 5574 38267
rect 14350 38233 14384 38267
rect 3985 38165 4019 38199
rect 10057 38165 10091 38199
rect 11989 38165 12023 38199
rect 13553 38165 13587 38199
rect 7389 37961 7423 37995
rect 12909 37961 12943 37995
rect 8125 37893 8159 37927
rect 2881 37825 2915 37859
rect 3893 37825 3927 37859
rect 4160 37825 4194 37859
rect 6837 37825 6871 37859
rect 6929 37825 6963 37859
rect 7113 37825 7147 37859
rect 7205 37825 7239 37859
rect 8217 37825 8251 37859
rect 8861 37825 8895 37859
rect 9597 37825 9631 37859
rect 9686 37831 9720 37865
rect 9786 37825 9820 37859
rect 9965 37825 9999 37859
rect 10609 37825 10643 37859
rect 11529 37825 11563 37859
rect 11796 37825 11830 37859
rect 14013 37825 14047 37859
rect 14197 37825 14231 37859
rect 3157 37757 3191 37791
rect 8769 37757 8803 37791
rect 10793 37757 10827 37791
rect 13829 37757 13863 37791
rect 2973 37621 3007 37655
rect 3065 37621 3099 37655
rect 5273 37621 5307 37655
rect 9321 37621 9355 37655
rect 10425 37621 10459 37655
rect 6653 37417 6687 37451
rect 7205 37417 7239 37451
rect 10425 37417 10459 37451
rect 11805 37417 11839 37451
rect 6561 37349 6595 37383
rect 10333 37349 10367 37383
rect 4997 37281 5031 37315
rect 8953 37281 8987 37315
rect 10241 37281 10275 37315
rect 12357 37281 12391 37315
rect 2237 37213 2271 37247
rect 2421 37213 2455 37247
rect 4077 37213 4111 37247
rect 4169 37213 4203 37247
rect 4261 37213 4295 37247
rect 4445 37213 4479 37247
rect 5089 37213 5123 37247
rect 6653 37213 6687 37247
rect 8125 37213 8159 37247
rect 9229 37213 9263 37247
rect 10517 37213 10551 37247
rect 11161 37213 11195 37247
rect 11345 37213 11379 37247
rect 11437 37213 11471 37247
rect 11529 37213 11563 37247
rect 12265 37213 12299 37247
rect 12449 37213 12483 37247
rect 2881 37145 2915 37179
rect 3065 37145 3099 37179
rect 3249 37145 3283 37179
rect 3801 37145 3835 37179
rect 6377 37145 6411 37179
rect 7297 37145 7331 37179
rect 7849 37145 7883 37179
rect 8033 37145 8067 37179
rect 2421 37077 2455 37111
rect 5457 37077 5491 37111
rect 7947 37077 7981 37111
rect 2881 36873 2915 36907
rect 4261 36873 4295 36907
rect 6561 36873 6595 36907
rect 7113 36873 7147 36907
rect 10517 36873 10551 36907
rect 13461 36873 13495 36907
rect 4721 36805 4755 36839
rect 5181 36805 5215 36839
rect 2513 36737 2547 36771
rect 3893 36737 3927 36771
rect 5089 36737 5123 36771
rect 5641 36737 5675 36771
rect 6653 36737 6687 36771
rect 8226 36737 8260 36771
rect 8493 36737 8527 36771
rect 9137 36737 9171 36771
rect 9404 36737 9438 36771
rect 13553 36737 13587 36771
rect 15577 36737 15611 36771
rect 2605 36669 2639 36703
rect 3801 36669 3835 36703
rect 4813 36669 4847 36703
rect 5733 36669 5767 36703
rect 15761 36669 15795 36703
rect 4905 36533 4939 36567
rect 15393 36533 15427 36567
rect 3893 36329 3927 36363
rect 4445 36329 4479 36363
rect 7849 36329 7883 36363
rect 10793 36329 10827 36363
rect 8217 36261 8251 36295
rect 16129 36261 16163 36295
rect 8953 36193 8987 36227
rect 3801 36125 3835 36159
rect 3985 36125 4019 36159
rect 4445 36125 4479 36159
rect 4629 36125 4663 36159
rect 8033 36125 8067 36159
rect 8309 36125 8343 36159
rect 10793 36125 10827 36159
rect 10977 36125 11011 36159
rect 14933 36125 14967 36159
rect 15117 36125 15151 36159
rect 9220 36057 9254 36091
rect 15853 36057 15887 36091
rect 10333 35989 10367 36023
rect 14749 35989 14783 36023
rect 15577 35989 15611 36023
rect 15761 35989 15795 36023
rect 15945 35989 15979 36023
rect 9137 35785 9171 35819
rect 14289 35785 14323 35819
rect 17141 35785 17175 35819
rect 14994 35717 15028 35751
rect 5089 35649 5123 35683
rect 9413 35649 9447 35683
rect 9505 35649 9539 35683
rect 9597 35649 9631 35683
rect 9781 35649 9815 35683
rect 14105 35649 14139 35683
rect 16681 35649 16715 35683
rect 16957 35649 16991 35683
rect 1409 35581 1443 35615
rect 1685 35581 1719 35615
rect 14749 35581 14783 35615
rect 16773 35581 16807 35615
rect 5181 35445 5215 35479
rect 16129 35445 16163 35479
rect 16681 35445 16715 35479
rect 16773 35241 16807 35275
rect 7941 35173 7975 35207
rect 15393 35105 15427 35139
rect 14381 35037 14415 35071
rect 14473 35037 14507 35071
rect 14703 35037 14737 35071
rect 14841 35037 14875 35071
rect 8125 34969 8159 35003
rect 14565 34969 14599 35003
rect 15660 34969 15694 35003
rect 14197 34901 14231 34935
rect 10425 34697 10459 34731
rect 16681 34697 16715 34731
rect 12541 34629 12575 34663
rect 14298 34629 14332 34663
rect 10517 34561 10551 34595
rect 11805 34561 11839 34595
rect 11989 34561 12023 34595
rect 14565 34561 14599 34595
rect 15301 34561 15335 34595
rect 16865 34561 16899 34595
rect 12725 34493 12759 34527
rect 15025 34493 15059 34527
rect 11989 34357 12023 34391
rect 13185 34357 13219 34391
rect 7849 34153 7883 34187
rect 14289 34153 14323 34187
rect 16037 34153 16071 34187
rect 15669 34017 15703 34051
rect 6009 33949 6043 33983
rect 6101 33949 6135 33983
rect 6561 33949 6595 33983
rect 6745 33949 6779 33983
rect 7941 33949 7975 33983
rect 13369 33949 13403 33983
rect 14105 33949 14139 33983
rect 15853 33949 15887 33983
rect 5825 33881 5859 33915
rect 13124 33881 13158 33915
rect 5923 33813 5957 33847
rect 6653 33813 6687 33847
rect 11989 33813 12023 33847
rect 10977 33609 11011 33643
rect 7573 33541 7607 33575
rect 8401 33541 8435 33575
rect 13185 33541 13219 33575
rect 4712 33473 4746 33507
rect 6377 33473 6411 33507
rect 6561 33473 6595 33507
rect 8125 33473 8159 33507
rect 8217 33473 8251 33507
rect 8861 33473 8895 33507
rect 10701 33473 10735 33507
rect 10793 33473 10827 33507
rect 11897 33473 11931 33507
rect 11989 33473 12023 33507
rect 12265 33473 12299 33507
rect 14749 33473 14783 33507
rect 4445 33405 4479 33439
rect 6837 33405 6871 33439
rect 9137 33405 9171 33439
rect 12725 33405 12759 33439
rect 15025 33405 15059 33439
rect 7389 33337 7423 33371
rect 8401 33337 8435 33371
rect 9045 33337 9079 33371
rect 12817 33337 12851 33371
rect 5825 33269 5859 33303
rect 6745 33269 6779 33303
rect 8953 33269 8987 33303
rect 11713 33269 11747 33303
rect 12173 33269 12207 33303
rect 8217 33065 8251 33099
rect 8401 33065 8435 33099
rect 11529 33065 11563 33099
rect 14105 33065 14139 33099
rect 10057 32997 10091 33031
rect 10793 32997 10827 33031
rect 3893 32929 3927 32963
rect 14473 32929 14507 32963
rect 15393 32929 15427 32963
rect 3985 32861 4019 32895
rect 4721 32861 4755 32895
rect 4997 32861 5031 32895
rect 5273 32861 5307 32895
rect 5549 32861 5583 32895
rect 6009 32861 6043 32895
rect 9137 32861 9171 32895
rect 9321 32861 9355 32895
rect 12909 32861 12943 32895
rect 14289 32861 14323 32895
rect 15117 32861 15151 32895
rect 3801 32793 3835 32827
rect 4261 32793 4295 32827
rect 6276 32793 6310 32827
rect 8033 32793 8067 32827
rect 8233 32793 8267 32827
rect 8953 32793 8987 32827
rect 10241 32793 10275 32827
rect 10977 32793 11011 32827
rect 12642 32793 12676 32827
rect 4169 32725 4203 32759
rect 4813 32725 4847 32759
rect 7389 32725 7423 32759
rect 6469 32521 6503 32555
rect 6637 32521 6671 32555
rect 7573 32521 7607 32555
rect 8861 32521 8895 32555
rect 10149 32521 10183 32555
rect 13185 32521 13219 32555
rect 6837 32453 6871 32487
rect 10057 32453 10091 32487
rect 10793 32453 10827 32487
rect 11713 32453 11747 32487
rect 13737 32453 13771 32487
rect 3617 32385 3651 32419
rect 3884 32385 3918 32419
rect 5641 32385 5675 32419
rect 5825 32385 5859 32419
rect 7298 32385 7332 32419
rect 8861 32385 8895 32419
rect 11897 32385 11931 32419
rect 11989 32385 12023 32419
rect 12265 32385 12299 32419
rect 7389 32317 7423 32351
rect 7573 32317 7607 32351
rect 8309 32317 8343 32351
rect 8953 32317 8987 32351
rect 12725 32317 12759 32351
rect 5825 32249 5859 32283
rect 12173 32249 12207 32283
rect 13093 32249 13127 32283
rect 4997 32181 5031 32215
rect 6653 32181 6687 32215
rect 10885 32181 10919 32215
rect 13829 32181 13863 32215
rect 4261 31977 4295 32011
rect 4813 31977 4847 32011
rect 5457 31977 5491 32011
rect 7757 31977 7791 32011
rect 9137 31977 9171 32011
rect 12725 31977 12759 32011
rect 7297 31909 7331 31943
rect 10977 31909 11011 31943
rect 3893 31841 3927 31875
rect 5825 31841 5859 31875
rect 9229 31841 9263 31875
rect 10149 31841 10183 31875
rect 11161 31841 11195 31875
rect 11713 31841 11747 31875
rect 3985 31773 4019 31807
rect 4813 31773 4847 31807
rect 4997 31773 5031 31807
rect 5641 31773 5675 31807
rect 5917 31773 5951 31807
rect 6009 31773 6043 31807
rect 6193 31773 6227 31807
rect 6653 31773 6687 31807
rect 6746 31773 6780 31807
rect 7021 31773 7055 31807
rect 7118 31773 7152 31807
rect 7941 31773 7975 31807
rect 8033 31773 8067 31807
rect 8953 31773 8987 31807
rect 9045 31773 9079 31807
rect 10057 31773 10091 31807
rect 10701 31773 10735 31807
rect 11897 31773 11931 31807
rect 12081 31773 12115 31807
rect 12541 31773 12575 31807
rect 6929 31705 6963 31739
rect 9689 31637 9723 31671
rect 10793 31637 10827 31671
rect 2881 31433 2915 31467
rect 5181 31433 5215 31467
rect 10333 31433 10367 31467
rect 11529 31365 11563 31399
rect 2513 31297 2547 31331
rect 3525 31297 3559 31331
rect 4353 31297 4387 31331
rect 5089 31297 5123 31331
rect 7021 31297 7055 31331
rect 8585 31297 8619 31331
rect 8677 31297 8711 31331
rect 8769 31297 8803 31331
rect 8953 31297 8987 31331
rect 9873 31297 9907 31331
rect 9965 31297 9999 31331
rect 10149 31297 10183 31331
rect 11805 31297 11839 31331
rect 14381 31297 14415 31331
rect 16865 31297 16899 31331
rect 2605 31229 2639 31263
rect 3341 31229 3375 31263
rect 4077 31229 4111 31263
rect 7297 31229 7331 31263
rect 11529 31229 11563 31263
rect 14565 31229 14599 31263
rect 10057 31161 10091 31195
rect 4169 31093 4203 31127
rect 4261 31093 4295 31127
rect 6837 31093 6871 31127
rect 7205 31093 7239 31127
rect 8309 31093 8343 31127
rect 11713 31093 11747 31127
rect 14197 31093 14231 31127
rect 16681 31093 16715 31127
rect 2697 30889 2731 30923
rect 4077 30889 4111 30923
rect 9045 30889 9079 30923
rect 10701 30889 10735 30923
rect 3065 30821 3099 30855
rect 10793 30753 10827 30787
rect 2881 30685 2915 30719
rect 2973 30685 3007 30719
rect 3157 30685 3191 30719
rect 3801 30685 3835 30719
rect 6469 30685 6503 30719
rect 8953 30685 8987 30719
rect 9137 30685 9171 30719
rect 10517 30685 10551 30719
rect 10609 30685 10643 30719
rect 13369 30685 13403 30719
rect 15485 30685 15519 30719
rect 17325 30685 17359 30719
rect 4077 30617 4111 30651
rect 6736 30617 6770 30651
rect 9689 30617 9723 30651
rect 9873 30617 9907 30651
rect 15240 30617 15274 30651
rect 17080 30617 17114 30651
rect 3893 30549 3927 30583
rect 7849 30549 7883 30583
rect 10057 30549 10091 30583
rect 13553 30549 13587 30583
rect 14105 30549 14139 30583
rect 15945 30549 15979 30583
rect 9137 30345 9171 30379
rect 15761 30345 15795 30379
rect 16681 30345 16715 30379
rect 17509 30345 17543 30379
rect 8024 30277 8058 30311
rect 7757 30209 7791 30243
rect 9873 30209 9907 30243
rect 10057 30209 10091 30243
rect 10517 30209 10551 30243
rect 10701 30209 10735 30243
rect 13921 30209 13955 30243
rect 14177 30209 14211 30243
rect 15945 30209 15979 30243
rect 16865 30209 16899 30243
rect 17693 30209 17727 30243
rect 9965 30141 9999 30175
rect 17049 30141 17083 30175
rect 10609 30005 10643 30039
rect 15301 30005 15335 30039
rect 5457 29801 5491 29835
rect 12725 29801 12759 29835
rect 14289 29801 14323 29835
rect 3249 29733 3283 29767
rect 13553 29733 13587 29767
rect 5825 29665 5859 29699
rect 9689 29665 9723 29699
rect 13185 29665 13219 29699
rect 16221 29665 16255 29699
rect 3065 29597 3099 29631
rect 3249 29597 3283 29631
rect 5641 29597 5675 29631
rect 5917 29597 5951 29631
rect 6009 29597 6043 29631
rect 6193 29597 6227 29631
rect 9597 29597 9631 29631
rect 11345 29597 11379 29631
rect 13369 29597 13403 29631
rect 14289 29597 14323 29631
rect 14381 29597 14415 29631
rect 15025 29597 15059 29631
rect 15209 29597 15243 29631
rect 11612 29529 11646 29563
rect 14565 29529 14599 29563
rect 16488 29529 16522 29563
rect 9965 29461 9999 29495
rect 14105 29461 14139 29495
rect 15393 29461 15427 29495
rect 17601 29461 17635 29495
rect 2881 29257 2915 29291
rect 5181 29257 5215 29291
rect 13829 29257 13863 29291
rect 15669 29257 15703 29291
rect 17049 29257 17083 29291
rect 14964 29189 14998 29223
rect 2513 29121 2547 29155
rect 3525 29121 3559 29155
rect 4169 29121 4203 29155
rect 5089 29121 5123 29155
rect 15209 29121 15243 29155
rect 15853 29121 15887 29155
rect 16773 29121 16807 29155
rect 16865 29121 16899 29155
rect 2605 29053 2639 29087
rect 3341 29053 3375 29087
rect 3709 29053 3743 29087
rect 4261 29053 4295 29087
rect 4445 29053 4479 29087
rect 4353 28917 4387 28951
rect 6285 28713 6319 28747
rect 12081 28713 12115 28747
rect 17141 28713 17175 28747
rect 14657 28645 14691 28679
rect 12449 28577 12483 28611
rect 13093 28577 13127 28611
rect 15761 28577 15795 28611
rect 3893 28509 3927 28543
rect 5733 28509 5767 28543
rect 6009 28509 6043 28543
rect 6101 28509 6135 28543
rect 7297 28509 7331 28543
rect 7481 28509 7515 28543
rect 10149 28509 10183 28543
rect 10333 28509 10367 28543
rect 12265 28509 12299 28543
rect 12357 28509 12391 28543
rect 12541 28509 12575 28543
rect 13277 28509 13311 28543
rect 14381 28509 14415 28543
rect 14473 28509 14507 28543
rect 4138 28441 4172 28475
rect 5917 28441 5951 28475
rect 14105 28441 14139 28475
rect 14289 28441 14323 28475
rect 16028 28441 16062 28475
rect 5273 28373 5307 28407
rect 7389 28373 7423 28407
rect 10241 28373 10275 28407
rect 13461 28373 13495 28407
rect 3801 28169 3835 28203
rect 7189 28169 7223 28203
rect 7849 28169 7883 28203
rect 12725 28169 12759 28203
rect 13185 28169 13219 28203
rect 16681 28169 16715 28203
rect 7389 28101 7423 28135
rect 4077 28033 4111 28067
rect 4169 28033 4203 28067
rect 4261 28033 4295 28067
rect 4445 28033 4479 28067
rect 8125 28033 8159 28067
rect 12081 28033 12115 28067
rect 12265 28033 12299 28067
rect 12357 28033 12391 28067
rect 12449 28033 12483 28067
rect 14298 28033 14332 28067
rect 14565 28033 14599 28067
rect 16865 28033 16899 28067
rect 7849 27965 7883 27999
rect 7021 27897 7055 27931
rect 7205 27829 7239 27863
rect 8033 27829 8067 27863
rect 5917 27625 5951 27659
rect 8309 27625 8343 27659
rect 13369 27625 13403 27659
rect 14289 27625 14323 27659
rect 10517 27557 10551 27591
rect 13553 27557 13587 27591
rect 6929 27421 6963 27455
rect 9689 27421 9723 27455
rect 9781 27421 9815 27455
rect 9873 27421 9907 27455
rect 10057 27421 10091 27455
rect 11345 27421 11379 27455
rect 11612 27421 11646 27455
rect 14105 27421 14139 27455
rect 5549 27353 5583 27387
rect 5733 27353 5767 27387
rect 7196 27353 7230 27387
rect 10701 27353 10735 27387
rect 13185 27353 13219 27387
rect 13401 27353 13435 27387
rect 9413 27285 9447 27319
rect 12725 27285 12759 27319
rect 5089 27081 5123 27115
rect 10517 27081 10551 27115
rect 11529 27081 11563 27115
rect 12173 27081 12207 27115
rect 17049 27081 17083 27115
rect 9404 27013 9438 27047
rect 12633 27013 12667 27047
rect 1685 26945 1719 26979
rect 4997 26945 5031 26979
rect 8410 26945 8444 26979
rect 8677 26945 8711 26979
rect 9137 26945 9171 26979
rect 11713 26945 11747 26979
rect 12357 26945 12391 26979
rect 16773 26945 16807 26979
rect 16865 26945 16899 26979
rect 12541 26877 12575 26911
rect 7297 26809 7331 26843
rect 1501 26741 1535 26775
rect 12449 26741 12483 26775
rect 4445 26537 4479 26571
rect 7757 26537 7791 26571
rect 8401 26537 8435 26571
rect 12081 26537 12115 26571
rect 11253 26469 11287 26503
rect 9873 26401 9907 26435
rect 12449 26401 12483 26435
rect 4583 26333 4617 26367
rect 4721 26333 4755 26367
rect 4996 26333 5030 26367
rect 5089 26333 5123 26367
rect 6929 26333 6963 26367
rect 7389 26333 7423 26367
rect 7573 26333 7607 26367
rect 8217 26333 8251 26367
rect 8401 26333 8435 26367
rect 9137 26333 9171 26367
rect 9229 26333 9263 26367
rect 12265 26333 12299 26367
rect 4813 26265 4847 26299
rect 6662 26265 6696 26299
rect 9413 26265 9447 26299
rect 10140 26265 10174 26299
rect 5549 26197 5583 26231
rect 6377 25993 6411 26027
rect 8033 25993 8067 26027
rect 9873 25993 9907 26027
rect 10517 25993 10551 26027
rect 11529 25993 11563 26027
rect 6653 25925 6687 25959
rect 3617 25857 3651 25891
rect 3873 25857 3907 25891
rect 6377 25857 6411 25891
rect 7757 25857 7791 25891
rect 9965 25857 9999 25891
rect 10701 25857 10735 25891
rect 12653 25857 12687 25891
rect 12909 25857 12943 25891
rect 15485 25857 15519 25891
rect 16681 25857 16715 25891
rect 7849 25789 7883 25823
rect 8033 25789 8067 25823
rect 16773 25789 16807 25823
rect 6469 25721 6503 25755
rect 4997 25653 5031 25687
rect 15669 25653 15703 25687
rect 16865 25653 16899 25687
rect 17049 25653 17083 25687
rect 3801 25449 3835 25483
rect 5273 25449 5307 25483
rect 6193 25449 6227 25483
rect 6377 25449 6411 25483
rect 13277 25449 13311 25483
rect 16589 25449 16623 25483
rect 11989 25313 12023 25347
rect 4077 25245 4111 25279
rect 4169 25245 4203 25279
rect 4261 25245 4295 25279
rect 4445 25245 4479 25279
rect 5273 25245 5307 25279
rect 5549 25245 5583 25279
rect 9689 25245 9723 25279
rect 9781 25245 9815 25279
rect 10977 25245 11011 25279
rect 11621 25245 11655 25279
rect 11805 25245 11839 25279
rect 12541 25245 12575 25279
rect 12633 25245 12667 25279
rect 12817 25245 12851 25279
rect 13461 25245 13495 25279
rect 14473 25245 14507 25279
rect 15485 25245 15519 25279
rect 15577 25245 15611 25279
rect 15945 25245 15979 25279
rect 6009 25177 6043 25211
rect 6209 25177 6243 25211
rect 9965 25177 9999 25211
rect 15669 25177 15703 25211
rect 15807 25177 15841 25211
rect 16773 25177 16807 25211
rect 5457 25109 5491 25143
rect 11161 25109 11195 25143
rect 14657 25109 14691 25143
rect 15301 25109 15335 25143
rect 16405 25109 16439 25143
rect 16573 25109 16607 25143
rect 12909 24905 12943 24939
rect 14289 24905 14323 24939
rect 11774 24837 11808 24871
rect 5089 24769 5123 24803
rect 5273 24769 5307 24803
rect 5457 24769 5491 24803
rect 5641 24769 5675 24803
rect 5825 24769 5859 24803
rect 14105 24769 14139 24803
rect 15016 24769 15050 24803
rect 16681 24769 16715 24803
rect 16865 24769 16899 24803
rect 16957 24769 16991 24803
rect 17141 24769 17175 24803
rect 17877 24769 17911 24803
rect 18153 24769 18187 24803
rect 5549 24701 5583 24735
rect 11529 24701 11563 24735
rect 13921 24701 13955 24735
rect 14749 24701 14783 24735
rect 17969 24701 18003 24735
rect 16129 24633 16163 24667
rect 17049 24633 17083 24667
rect 17693 24633 17727 24667
rect 17877 24565 17911 24599
rect 5181 24361 5215 24395
rect 14749 24361 14783 24395
rect 16589 24361 16623 24395
rect 17141 24361 17175 24395
rect 2513 24225 2547 24259
rect 3801 24225 3835 24259
rect 3985 24225 4019 24259
rect 14381 24225 14415 24259
rect 2605 24157 2639 24191
rect 4077 24157 4111 24191
rect 5273 24157 5307 24191
rect 14565 24157 14599 24191
rect 15209 24157 15243 24191
rect 17325 24157 17359 24191
rect 12449 24089 12483 24123
rect 15476 24089 15510 24123
rect 17509 24089 17543 24123
rect 17693 24089 17727 24123
rect 2973 24021 3007 24055
rect 3801 24021 3835 24055
rect 11161 24021 11195 24055
rect 17417 24021 17451 24055
rect 3249 23817 3283 23851
rect 18153 23817 18187 23851
rect 3893 23749 3927 23783
rect 2973 23681 3007 23715
rect 3157 23681 3191 23715
rect 4077 23681 4111 23715
rect 7205 23681 7239 23715
rect 7665 23681 7699 23715
rect 7849 23681 7883 23715
rect 13093 23681 13127 23715
rect 13277 23681 13311 23715
rect 14850 23681 14884 23715
rect 15117 23681 15151 23715
rect 16129 23681 16163 23715
rect 16773 23681 16807 23715
rect 17040 23681 17074 23715
rect 3433 23477 3467 23511
rect 7021 23477 7055 23511
rect 7849 23477 7883 23511
rect 13277 23477 13311 23511
rect 13737 23477 13771 23511
rect 15945 23477 15979 23511
rect 2697 23273 2731 23307
rect 3801 23273 3835 23307
rect 5549 23273 5583 23307
rect 9137 23273 9171 23307
rect 3065 23205 3099 23239
rect 6101 23205 6135 23239
rect 8953 23205 8987 23239
rect 14289 23205 14323 23239
rect 3985 23137 4019 23171
rect 4077 23137 4111 23171
rect 13461 23137 13495 23171
rect 14105 23137 14139 23171
rect 15393 23137 15427 23171
rect 15945 23137 15979 23171
rect 16773 23137 16807 23171
rect 2881 23069 2915 23103
rect 2973 23069 3007 23103
rect 3157 23069 3191 23103
rect 5365 23069 5399 23103
rect 5641 23069 5675 23103
rect 6377 23069 6411 23103
rect 7021 23069 7055 23103
rect 8309 23069 8343 23103
rect 8401 23069 8435 23103
rect 13185 23069 13219 23103
rect 13277 23069 13311 23103
rect 13553 23069 13587 23103
rect 15209 23069 15243 23103
rect 16129 23069 16163 23103
rect 6101 23001 6135 23035
rect 7389 23001 7423 23035
rect 8125 23001 8159 23035
rect 9105 23001 9139 23035
rect 9321 23001 9355 23035
rect 14565 23001 14599 23035
rect 17040 23001 17074 23035
rect 4445 22933 4479 22967
rect 5181 22933 5215 22967
rect 6285 22933 6319 22967
rect 8401 22933 8435 22967
rect 13001 22933 13035 22967
rect 15025 22933 15059 22967
rect 16313 22933 16347 22967
rect 18153 22933 18187 22967
rect 3249 22729 3283 22763
rect 3801 22729 3835 22763
rect 10339 22729 10373 22763
rect 14105 22729 14139 22763
rect 3893 22661 3927 22695
rect 8646 22661 8680 22695
rect 10425 22661 10459 22695
rect 2973 22593 3007 22627
rect 4445 22593 4479 22627
rect 4712 22593 4746 22627
rect 6929 22593 6963 22627
rect 10241 22593 10275 22627
rect 10517 22593 10551 22627
rect 11529 22593 11563 22627
rect 12532 22593 12566 22627
rect 15025 22593 15059 22627
rect 15301 22593 15335 22627
rect 16681 22593 16715 22627
rect 16948 22593 16982 22627
rect 3249 22525 3283 22559
rect 7205 22525 7239 22559
rect 8401 22525 8435 22559
rect 12265 22525 12299 22559
rect 14565 22525 14599 22559
rect 3065 22457 3099 22491
rect 13645 22457 13679 22491
rect 14289 22457 14323 22491
rect 5825 22389 5859 22423
rect 9781 22389 9815 22423
rect 11713 22389 11747 22423
rect 18061 22389 18095 22423
rect 3157 22185 3191 22219
rect 13461 22185 13495 22219
rect 3893 22049 3927 22083
rect 5733 22049 5767 22083
rect 6009 22049 6043 22083
rect 9597 22049 9631 22083
rect 13553 22049 13587 22083
rect 17969 22049 18003 22083
rect 2421 21981 2455 22015
rect 2605 21981 2639 22015
rect 3065 21981 3099 22015
rect 3249 21981 3283 22015
rect 4077 21981 4111 22015
rect 5273 21981 5307 22015
rect 7021 21981 7055 22015
rect 9137 21981 9171 22015
rect 11437 21981 11471 22015
rect 11621 21981 11655 22015
rect 13185 21981 13219 22015
rect 13277 21981 13311 22015
rect 14473 21981 14507 22015
rect 14565 21981 14599 22015
rect 16129 21981 16163 22015
rect 16773 21981 16807 22015
rect 16957 21981 16991 22015
rect 17141 21981 17175 22015
rect 17785 21981 17819 22015
rect 4261 21913 4295 21947
rect 7288 21913 7322 21947
rect 9864 21913 9898 21947
rect 11529 21913 11563 21947
rect 13001 21913 13035 21947
rect 2605 21845 2639 21879
rect 5089 21845 5123 21879
rect 8401 21845 8435 21879
rect 9045 21845 9079 21879
rect 10977 21845 11011 21879
rect 14289 21845 14323 21879
rect 16313 21845 16347 21879
rect 17601 21845 17635 21879
rect 5825 21641 5859 21675
rect 10425 21641 10459 21675
rect 13277 21641 13311 21675
rect 17141 21641 17175 21675
rect 17601 21641 17635 21675
rect 2881 21505 2915 21539
rect 4077 21505 4111 21539
rect 4169 21505 4203 21539
rect 4261 21505 4295 21539
rect 4445 21505 4479 21539
rect 5273 21505 5307 21539
rect 5365 21505 5399 21539
rect 5549 21505 5583 21539
rect 5641 21505 5675 21539
rect 7490 21505 7524 21539
rect 7757 21505 7791 21539
rect 8217 21505 8251 21539
rect 8484 21505 8518 21539
rect 10241 21505 10275 21539
rect 11529 21505 11563 21539
rect 13461 21505 13495 21539
rect 16957 21505 16991 21539
rect 17785 21505 17819 21539
rect 2789 21437 2823 21471
rect 10057 21437 10091 21471
rect 3249 21369 3283 21403
rect 6377 21369 6411 21403
rect 3801 21301 3835 21335
rect 9597 21301 9631 21335
rect 11713 21301 11747 21335
rect 5273 21097 5307 21131
rect 17877 21097 17911 21131
rect 6193 20961 6227 20995
rect 6469 20961 6503 20995
rect 11345 20961 11379 20995
rect 3893 20893 3927 20927
rect 7849 20893 7883 20927
rect 8125 20893 8159 20927
rect 10885 20893 10919 20927
rect 11612 20893 11646 20927
rect 13277 20893 13311 20927
rect 13369 20893 13403 20927
rect 18061 20893 18095 20927
rect 4138 20825 4172 20859
rect 8033 20825 8067 20859
rect 10640 20825 10674 20859
rect 7665 20757 7699 20791
rect 9505 20757 9539 20791
rect 12725 20757 12759 20791
rect 3893 20553 3927 20587
rect 5733 20553 5767 20587
rect 7757 20553 7791 20587
rect 10083 20553 10117 20587
rect 10977 20553 11011 20587
rect 7573 20485 7607 20519
rect 9873 20485 9907 20519
rect 11989 20485 12023 20519
rect 13093 20485 13127 20519
rect 3709 20417 3743 20451
rect 3893 20417 3927 20451
rect 5641 20417 5675 20451
rect 5825 20417 5859 20451
rect 6653 20417 6687 20451
rect 7849 20417 7883 20451
rect 9045 20417 9079 20451
rect 10701 20417 10735 20451
rect 10793 20417 10827 20451
rect 12909 20417 12943 20451
rect 10977 20349 11011 20383
rect 7573 20281 7607 20315
rect 12173 20281 12207 20315
rect 6469 20213 6503 20247
rect 8953 20213 8987 20247
rect 10057 20213 10091 20247
rect 10241 20213 10275 20247
rect 8125 20009 8159 20043
rect 10793 20009 10827 20043
rect 10149 19941 10183 19975
rect 14749 19941 14783 19975
rect 10333 19873 10367 19907
rect 8217 19805 8251 19839
rect 9597 19805 9631 19839
rect 10057 19805 10091 19839
rect 10793 19805 10827 19839
rect 10977 19805 11011 19839
rect 15577 19805 15611 19839
rect 15761 19805 15795 19839
rect 10333 19737 10367 19771
rect 14565 19737 14599 19771
rect 9505 19669 9539 19703
rect 15945 19669 15979 19703
rect 14749 19465 14783 19499
rect 9505 19397 9539 19431
rect 14289 19397 14323 19431
rect 9597 19329 9631 19363
rect 12909 19329 12943 19363
rect 14473 19329 14507 19363
rect 14565 19329 14599 19363
rect 16681 19329 16715 19363
rect 13093 19261 13127 19295
rect 15209 19261 15243 19295
rect 15485 19261 15519 19295
rect 14289 19125 14323 19159
rect 16865 19125 16899 19159
rect 5641 18921 5675 18955
rect 14381 18921 14415 18955
rect 16221 18921 16255 18955
rect 12449 18853 12483 18887
rect 13185 18785 13219 18819
rect 5733 18717 5767 18751
rect 12265 18717 12299 18751
rect 12449 18717 12483 18751
rect 13369 18717 13403 18751
rect 15761 18717 15795 18751
rect 17601 18717 17635 18751
rect 15494 18649 15528 18683
rect 17334 18649 17368 18683
rect 13553 18581 13587 18615
rect 4905 18377 4939 18411
rect 7481 18309 7515 18343
rect 4813 18241 4847 18275
rect 5733 18241 5767 18275
rect 6469 18241 6503 18275
rect 6561 18241 6595 18275
rect 6745 18241 6779 18275
rect 7205 18241 7239 18275
rect 12449 18241 12483 18275
rect 14666 18241 14700 18275
rect 14933 18241 14967 18275
rect 15393 18241 15427 18275
rect 15577 18241 15611 18275
rect 15669 18241 15703 18275
rect 15761 18241 15795 18275
rect 16865 18241 16899 18275
rect 7481 18173 7515 18207
rect 12633 18173 12667 18207
rect 17049 18173 17083 18207
rect 6745 18105 6779 18139
rect 1409 18037 1443 18071
rect 5549 18037 5583 18071
rect 7297 18037 7331 18071
rect 12265 18037 12299 18071
rect 13553 18037 13587 18071
rect 16037 18037 16071 18071
rect 16681 18037 16715 18071
rect 4997 17833 5031 17867
rect 7205 17833 7239 17867
rect 10793 17833 10827 17867
rect 16129 17833 16163 17867
rect 4445 17765 4479 17799
rect 11989 17765 12023 17799
rect 15485 17765 15519 17799
rect 6193 17697 6227 17731
rect 8033 17697 8067 17731
rect 12081 17697 12115 17731
rect 4261 17629 4295 17663
rect 5181 17629 5215 17663
rect 6285 17629 6319 17663
rect 6469 17629 6503 17663
rect 8217 17629 8251 17663
rect 9781 17629 9815 17663
rect 9965 17629 9999 17663
rect 11713 17629 11747 17663
rect 11805 17629 11839 17663
rect 12725 17629 12759 17663
rect 12817 17629 12851 17663
rect 13369 17629 13403 17663
rect 14105 17629 14139 17663
rect 16773 17629 16807 17663
rect 16957 17629 16991 17663
rect 17141 17629 17175 17663
rect 17785 17629 17819 17663
rect 7389 17561 7423 17595
rect 7573 17561 7607 17595
rect 10885 17561 10919 17595
rect 14350 17561 14384 17595
rect 16313 17561 16347 17595
rect 6653 17493 6687 17527
rect 9873 17493 9907 17527
rect 11529 17493 11563 17527
rect 12541 17493 12575 17527
rect 13553 17493 13587 17527
rect 15945 17493 15979 17527
rect 16113 17493 16147 17527
rect 17601 17493 17635 17527
rect 11621 17289 11655 17323
rect 14565 17289 14599 17323
rect 15577 17289 15611 17323
rect 18061 17289 18095 17323
rect 6644 17221 6678 17255
rect 10793 17221 10827 17255
rect 4169 17153 4203 17187
rect 4261 17153 4295 17187
rect 4353 17156 4387 17190
rect 4537 17153 4571 17187
rect 5181 17153 5215 17187
rect 5365 17153 5399 17187
rect 8217 17153 8251 17187
rect 8401 17153 8435 17187
rect 8585 17153 8619 17187
rect 8769 17153 8803 17187
rect 9873 17153 9907 17187
rect 10057 17153 10091 17187
rect 11805 17153 11839 17187
rect 11897 17153 11931 17187
rect 12173 17153 12207 17187
rect 13737 17153 13771 17187
rect 14841 17153 14875 17187
rect 15025 17153 15059 17187
rect 15761 17153 15795 17187
rect 16681 17153 16715 17187
rect 16948 17153 16982 17187
rect 5457 17085 5491 17119
rect 6377 17085 6411 17119
rect 8493 17085 8527 17119
rect 10149 17085 10183 17119
rect 12633 17085 12667 17119
rect 13093 17085 13127 17119
rect 13553 17085 13587 17119
rect 14749 17085 14783 17119
rect 14933 17085 14967 17119
rect 10977 17017 11011 17051
rect 12725 17017 12759 17051
rect 3893 16949 3927 16983
rect 4997 16949 5031 16983
rect 7757 16949 7791 16983
rect 8953 16949 8987 16983
rect 9689 16949 9723 16983
rect 12081 16949 12115 16983
rect 13921 16949 13955 16983
rect 3249 16745 3283 16779
rect 10701 16745 10735 16779
rect 14197 16745 14231 16779
rect 13093 16677 13127 16711
rect 13277 16677 13311 16711
rect 7021 16609 7055 16643
rect 9321 16609 9355 16643
rect 11253 16609 11287 16643
rect 13553 16609 13587 16643
rect 17417 16609 17451 16643
rect 2973 16541 3007 16575
rect 4077 16541 4111 16575
rect 4344 16541 4378 16575
rect 6193 16541 6227 16575
rect 6285 16541 6319 16575
rect 6377 16541 6411 16575
rect 6561 16541 6595 16575
rect 15025 16541 15059 16575
rect 17161 16541 17195 16575
rect 3249 16473 3283 16507
rect 5917 16473 5951 16507
rect 7266 16473 7300 16507
rect 9588 16473 9622 16507
rect 11520 16473 11554 16507
rect 14289 16473 14323 16507
rect 3065 16405 3099 16439
rect 5457 16405 5491 16439
rect 8401 16405 8435 16439
rect 12633 16405 12667 16439
rect 14841 16405 14875 16439
rect 16037 16405 16071 16439
rect 3709 16201 3743 16235
rect 6745 16201 6779 16235
rect 10977 16201 11011 16235
rect 11989 16201 12023 16235
rect 17325 16201 17359 16235
rect 2605 16133 2639 16167
rect 2805 16133 2839 16167
rect 6377 16133 6411 16167
rect 6593 16133 6627 16167
rect 9873 16133 9907 16167
rect 9965 16133 9999 16167
rect 3985 16065 4019 16099
rect 5549 16065 5583 16099
rect 5825 16065 5859 16099
rect 7757 16065 7791 16099
rect 8033 16065 8067 16099
rect 8493 16065 8527 16099
rect 8677 16065 8711 16099
rect 8953 16065 8987 16099
rect 9781 16065 9815 16099
rect 10149 16065 10183 16099
rect 10701 16065 10735 16099
rect 10793 16065 10827 16099
rect 13113 16065 13147 16099
rect 13369 16065 13403 16099
rect 17509 16065 17543 16099
rect 3433 15997 3467 16031
rect 4077 15997 4111 16031
rect 2789 15861 2823 15895
rect 2973 15861 3007 15895
rect 6561 15861 6595 15895
rect 9137 15861 9171 15895
rect 9597 15861 9631 15895
rect 5273 15657 5307 15691
rect 6101 15657 6135 15691
rect 7757 15657 7791 15691
rect 11529 15657 11563 15691
rect 3249 15589 3283 15623
rect 3893 15521 3927 15555
rect 6561 15521 6595 15555
rect 7205 15521 7239 15555
rect 10977 15521 11011 15555
rect 11713 15521 11747 15555
rect 2973 15453 3007 15487
rect 5825 15453 5859 15487
rect 5917 15453 5951 15487
rect 7113 15453 7147 15487
rect 7936 15453 7970 15487
rect 8253 15453 8287 15487
rect 8401 15453 8435 15487
rect 11437 15453 11471 15487
rect 12357 15453 12391 15487
rect 3249 15385 3283 15419
rect 4160 15385 4194 15419
rect 6101 15385 6135 15419
rect 8033 15385 8067 15419
rect 8125 15385 8159 15419
rect 10732 15385 10766 15419
rect 14197 15385 14231 15419
rect 14381 15385 14415 15419
rect 3065 15317 3099 15351
rect 6837 15317 6871 15351
rect 9597 15317 9631 15351
rect 11713 15317 11747 15351
rect 12173 15317 12207 15351
rect 3617 15113 3651 15147
rect 4077 15113 4111 15147
rect 7573 15113 7607 15147
rect 10133 15113 10167 15147
rect 10885 15113 10919 15147
rect 17509 15113 17543 15147
rect 4261 15045 4295 15079
rect 10333 15045 10367 15079
rect 11989 15045 12023 15079
rect 3341 14977 3375 15011
rect 3433 14977 3467 15011
rect 4445 14977 4479 15011
rect 6929 14977 6963 15011
rect 7573 14977 7607 15011
rect 7757 14977 7791 15011
rect 8585 14977 8619 15011
rect 8861 14977 8895 15011
rect 8953 14977 8987 15011
rect 10793 14977 10827 15011
rect 10977 14977 11011 15011
rect 17693 14977 17727 15011
rect 3617 14909 3651 14943
rect 8677 14909 8711 14943
rect 17877 14909 17911 14943
rect 7113 14841 7147 14875
rect 9965 14841 9999 14875
rect 9137 14773 9171 14807
rect 10149 14773 10183 14807
rect 12081 14773 12115 14807
rect 4077 14569 4111 14603
rect 9321 14569 9355 14603
rect 17969 14569 18003 14603
rect 9413 14433 9447 14467
rect 3985 14365 4019 14399
rect 4169 14365 4203 14399
rect 9137 14365 9171 14399
rect 10609 14365 10643 14399
rect 15761 14365 15795 14399
rect 18153 14365 18187 14399
rect 9873 14297 9907 14331
rect 10057 14297 10091 14331
rect 8953 14229 8987 14263
rect 10701 14229 10735 14263
rect 15577 14229 15611 14263
rect 15577 14025 15611 14059
rect 9597 13957 9631 13991
rect 9781 13957 9815 13991
rect 14565 13957 14599 13991
rect 13829 13889 13863 13923
rect 15761 13889 15795 13923
rect 13645 13821 13679 13855
rect 14013 13821 14047 13855
rect 15945 13821 15979 13855
rect 14749 13753 14783 13787
rect 15945 13481 15979 13515
rect 16957 13481 16991 13515
rect 17417 13481 17451 13515
rect 17049 13345 17083 13379
rect 13277 13277 13311 13311
rect 13369 13277 13403 13311
rect 15485 13277 15519 13311
rect 16313 13277 16347 13311
rect 16497 13277 16531 13311
rect 17233 13277 17267 13311
rect 15218 13209 15252 13243
rect 16129 13209 16163 13243
rect 16957 13209 16991 13243
rect 13553 13141 13587 13175
rect 14105 13141 14139 13175
rect 16221 13141 16255 13175
rect 13001 12937 13035 12971
rect 8585 12869 8619 12903
rect 9597 12869 9631 12903
rect 16129 12869 16163 12903
rect 10333 12801 10367 12835
rect 11888 12801 11922 12835
rect 14574 12801 14608 12835
rect 14841 12801 14875 12835
rect 15945 12801 15979 12835
rect 16865 12801 16899 12835
rect 17693 12801 17727 12835
rect 11621 12733 11655 12767
rect 15761 12733 15795 12767
rect 16681 12733 16715 12767
rect 8677 12597 8711 12631
rect 9505 12597 9539 12631
rect 10241 12597 10275 12631
rect 13461 12597 13495 12631
rect 17049 12597 17083 12631
rect 17509 12597 17543 12631
rect 8401 12393 8435 12427
rect 12357 12393 12391 12427
rect 14105 12393 14139 12427
rect 16773 12393 16807 12427
rect 10057 12325 10091 12359
rect 13553 12325 13587 12359
rect 10977 12257 11011 12291
rect 15393 12257 15427 12291
rect 7021 12189 7055 12223
rect 8953 12189 8987 12223
rect 9101 12189 9135 12223
rect 9229 12189 9263 12223
rect 9459 12189 9493 12223
rect 10333 12189 10367 12223
rect 13277 12189 13311 12223
rect 14289 12189 14323 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 14749 12189 14783 12223
rect 17417 12189 17451 12223
rect 7288 12121 7322 12155
rect 9321 12121 9355 12155
rect 10057 12121 10091 12155
rect 11244 12121 11278 12155
rect 13001 12121 13035 12155
rect 14591 12121 14625 12155
rect 15660 12121 15694 12155
rect 9597 12053 9631 12087
rect 10241 12053 10275 12087
rect 13185 12053 13219 12087
rect 13369 12053 13403 12087
rect 17233 12053 17267 12087
rect 6929 11849 6963 11883
rect 13921 11849 13955 11883
rect 16129 11849 16163 11883
rect 5825 11781 5859 11815
rect 9873 11781 9907 11815
rect 10793 11781 10827 11815
rect 15016 11781 15050 11815
rect 4905 11713 4939 11747
rect 5089 11713 5123 11747
rect 5549 11713 5583 11747
rect 5641 11713 5675 11747
rect 7205 11713 7239 11747
rect 7297 11713 7331 11747
rect 7389 11713 7423 11747
rect 7573 11713 7607 11747
rect 8861 11713 8895 11747
rect 9597 11713 9631 11747
rect 9690 11713 9724 11747
rect 9965 11713 9999 11747
rect 10103 11713 10137 11747
rect 10701 11713 10735 11747
rect 12081 11713 12115 11747
rect 12348 11713 12382 11747
rect 14105 11713 14139 11747
rect 14289 11713 14323 11747
rect 9137 11645 9171 11679
rect 14749 11645 14783 11679
rect 9045 11577 9079 11611
rect 4905 11509 4939 11543
rect 5825 11509 5859 11543
rect 8677 11509 8711 11543
rect 10241 11509 10275 11543
rect 13461 11509 13495 11543
rect 7757 11305 7791 11339
rect 10517 11305 10551 11339
rect 11529 11305 11563 11339
rect 14105 11305 14139 11339
rect 14565 11305 14599 11339
rect 15301 11305 15335 11339
rect 11713 11237 11747 11271
rect 6285 11169 6319 11203
rect 7665 11169 7699 11203
rect 9137 11169 9171 11203
rect 12173 11169 12207 11203
rect 12449 11169 12483 11203
rect 14197 11169 14231 11203
rect 3985 11101 4019 11135
rect 6193 11101 6227 11135
rect 6837 11101 6871 11135
rect 7021 11101 7055 11135
rect 7205 11101 7239 11135
rect 7849 11101 7883 11135
rect 7941 11101 7975 11135
rect 9393 11101 9427 11135
rect 14381 11101 14415 11135
rect 16681 11101 16715 11135
rect 4252 11033 4286 11067
rect 11345 11033 11379 11067
rect 14105 11033 14139 11067
rect 16436 11033 16470 11067
rect 5365 10965 5399 10999
rect 5825 10965 5859 10999
rect 11545 10965 11579 10999
rect 5181 10761 5215 10795
rect 8401 10761 8435 10795
rect 8953 10761 8987 10795
rect 10609 10761 10643 10795
rect 14013 10761 14047 10795
rect 14657 10761 14691 10795
rect 4261 10693 4295 10727
rect 4721 10693 4755 10727
rect 7665 10693 7699 10727
rect 12173 10693 12207 10727
rect 4445 10625 4479 10659
rect 4629 10625 4663 10659
rect 5549 10625 5583 10659
rect 6561 10625 6595 10659
rect 8309 10625 8343 10659
rect 8493 10625 8527 10659
rect 9137 10625 9171 10659
rect 9413 10625 9447 10659
rect 9505 10625 9539 10659
rect 9689 10625 9723 10659
rect 10149 10625 10183 10659
rect 13185 10625 13219 10659
rect 13829 10625 13863 10659
rect 14473 10625 14507 10659
rect 4353 10557 4387 10591
rect 5641 10557 5675 10591
rect 6469 10557 6503 10591
rect 9321 10557 9355 10591
rect 12449 10557 12483 10591
rect 13369 10557 13403 10591
rect 6929 10489 6963 10523
rect 7757 10421 7791 10455
rect 10425 10421 10459 10455
rect 13001 10421 13035 10455
rect 5181 10217 5215 10251
rect 11897 10217 11931 10251
rect 12725 10217 12759 10251
rect 6009 10149 6043 10183
rect 6101 10149 6135 10183
rect 6929 10149 6963 10183
rect 5365 10081 5399 10115
rect 6837 10081 6871 10115
rect 7849 10081 7883 10115
rect 11529 10081 11563 10115
rect 5089 10013 5123 10047
rect 5917 10013 5951 10047
rect 6193 10013 6227 10047
rect 7021 10013 7055 10047
rect 7113 10013 7147 10047
rect 7941 10013 7975 10047
rect 11437 10013 11471 10047
rect 11621 10013 11655 10047
rect 11713 10013 11747 10047
rect 12909 10013 12943 10047
rect 5365 9945 5399 9979
rect 6377 9877 6411 9911
rect 7573 9877 7607 9911
rect 6469 9605 6503 9639
rect 6653 9605 6687 9639
rect 7757 9605 7791 9639
rect 4997 9537 5031 9571
rect 5181 9537 5215 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 7573 9537 7607 9571
rect 9597 9537 9631 9571
rect 9864 9537 9898 9571
rect 7481 9401 7515 9435
rect 4997 9333 5031 9367
rect 10977 9333 11011 9367
rect 4721 9129 4755 9163
rect 10241 9129 10275 9163
rect 11161 9129 11195 9163
rect 7573 9061 7607 9095
rect 4629 8993 4663 9027
rect 11437 8993 11471 9027
rect 1409 8925 1443 8959
rect 4813 8925 4847 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 7389 8925 7423 8959
rect 10425 8925 10459 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 11657 8925 11691 8959
rect 4537 8857 4571 8891
rect 4997 8857 5031 8891
rect 5273 8585 5307 8619
rect 10425 8585 10459 8619
rect 12081 8585 12115 8619
rect 4160 8517 4194 8551
rect 11713 8517 11747 8551
rect 3893 8449 3927 8483
rect 7757 8449 7791 8483
rect 10609 8449 10643 8483
rect 11805 8449 11839 8483
rect 11897 8449 11931 8483
rect 14289 8449 14323 8483
rect 8033 8381 8067 8415
rect 10793 8381 10827 8415
rect 14473 8381 14507 8415
rect 7941 8313 7975 8347
rect 11529 8313 11563 8347
rect 7849 8245 7883 8279
rect 14105 8245 14139 8279
rect 8033 8041 8067 8075
rect 14565 8041 14599 8075
rect 14933 8041 14967 8075
rect 8217 7905 8251 7939
rect 14933 7905 14967 7939
rect 7757 7837 7791 7871
rect 7849 7837 7883 7871
rect 11805 7837 11839 7871
rect 12633 7837 12667 7871
rect 13369 7837 13403 7871
rect 14749 7837 14783 7871
rect 15025 7769 15059 7803
rect 11621 7701 11655 7735
rect 12817 7701 12851 7735
rect 13553 7701 13587 7735
rect 9505 7497 9539 7531
rect 11529 7497 11563 7531
rect 14258 7429 14292 7463
rect 8125 7361 8159 7395
rect 8392 7361 8426 7395
rect 10517 7361 10551 7395
rect 10701 7361 10735 7395
rect 11897 7361 11931 7395
rect 12633 7361 12667 7395
rect 11805 7293 11839 7327
rect 14013 7293 14047 7327
rect 10333 7157 10367 7191
rect 11897 7157 11931 7191
rect 12449 7157 12483 7191
rect 15393 7157 15427 7191
rect 8309 6953 8343 6987
rect 14933 6885 14967 6919
rect 15761 6885 15795 6919
rect 11897 6817 11931 6851
rect 14381 6817 14415 6851
rect 7665 6749 7699 6783
rect 7849 6749 7883 6783
rect 7941 6749 7975 6783
rect 8033 6749 8067 6783
rect 10241 6749 10275 6783
rect 12164 6749 12198 6783
rect 17141 6749 17175 6783
rect 14749 6681 14783 6715
rect 16874 6681 16908 6715
rect 10057 6613 10091 6647
rect 13277 6613 13311 6647
rect 14565 6613 14599 6647
rect 14657 6613 14691 6647
rect 7849 6409 7883 6443
rect 12173 6409 12207 6443
rect 12449 6409 12483 6443
rect 13185 6409 13219 6443
rect 14013 6409 14047 6443
rect 4905 6273 4939 6307
rect 6929 6273 6963 6307
rect 7113 6273 7147 6307
rect 7573 6273 7607 6307
rect 7665 6273 7699 6307
rect 12357 6273 12391 6307
rect 12541 6273 12575 6307
rect 13369 6273 13403 6307
rect 13461 6273 13495 6307
rect 15137 6273 15171 6307
rect 15393 6273 15427 6307
rect 16037 6273 16071 6307
rect 17325 6273 17359 6307
rect 17509 6273 17543 6307
rect 4997 6205 5031 6239
rect 7849 6205 7883 6239
rect 12725 6137 12759 6171
rect 15853 6137 15887 6171
rect 4537 6069 4571 6103
rect 7021 6069 7055 6103
rect 17141 6069 17175 6103
rect 4813 5865 4847 5899
rect 6745 5865 6779 5899
rect 10885 5865 10919 5899
rect 12173 5865 12207 5899
rect 12633 5865 12667 5899
rect 15485 5865 15519 5899
rect 16773 5865 16807 5899
rect 17969 5865 18003 5899
rect 4997 5729 5031 5763
rect 7113 5729 7147 5763
rect 9505 5729 9539 5763
rect 11345 5729 11379 5763
rect 12449 5729 12483 5763
rect 15117 5729 15151 5763
rect 5089 5661 5123 5695
rect 5917 5661 5951 5695
rect 6101 5661 6135 5695
rect 7021 5661 7055 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 9772 5661 9806 5695
rect 11529 5661 11563 5695
rect 12357 5661 12391 5695
rect 13093 5661 13127 5695
rect 13277 5661 13311 5695
rect 14381 5661 14415 5695
rect 14473 5661 14507 5695
rect 15301 5661 15335 5695
rect 16129 5661 16163 5695
rect 16221 5661 16255 5695
rect 16957 5661 16991 5695
rect 18153 5661 18187 5695
rect 11713 5593 11747 5627
rect 12633 5593 12667 5627
rect 6009 5525 6043 5559
rect 8125 5525 8159 5559
rect 13461 5525 13495 5559
rect 14657 5525 14691 5559
rect 15945 5525 15979 5559
rect 5273 5321 5307 5355
rect 12173 5321 12207 5355
rect 15393 5321 15427 5355
rect 6377 5253 6411 5287
rect 6745 5253 6779 5287
rect 8769 5253 8803 5287
rect 4629 5185 4663 5219
rect 4813 5185 4847 5219
rect 5549 5185 5583 5219
rect 6561 5185 6595 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 7573 5185 7607 5219
rect 7665 5185 7699 5219
rect 8585 5185 8619 5219
rect 9965 5185 9999 5219
rect 10425 5185 10459 5219
rect 10609 5185 10643 5219
rect 10793 5185 10827 5219
rect 11529 5185 11563 5219
rect 13297 5185 13331 5219
rect 13553 5185 13587 5219
rect 14013 5185 14047 5219
rect 14280 5185 14314 5219
rect 5273 5117 5307 5151
rect 4721 5049 4755 5083
rect 5457 4981 5491 5015
rect 7941 4981 7975 5015
rect 8401 4981 8435 5015
rect 9781 4981 9815 5015
rect 11713 4981 11747 5015
rect 7573 4777 7607 4811
rect 8217 4777 8251 4811
rect 10977 4777 11011 4811
rect 12817 4777 12851 4811
rect 14105 4777 14139 4811
rect 14749 4777 14783 4811
rect 5457 4641 5491 4675
rect 9597 4641 9631 4675
rect 11437 4641 11471 4675
rect 5365 4573 5399 4607
rect 6469 4573 6503 4607
rect 6558 4570 6592 4604
rect 6653 4573 6687 4607
rect 6837 4573 6871 4607
rect 7481 4573 7515 4607
rect 7665 4573 7699 4607
rect 9853 4573 9887 4607
rect 11704 4573 11738 4607
rect 13461 4573 13495 4607
rect 14289 4573 14323 4607
rect 14933 4573 14967 4607
rect 15577 4573 15611 4607
rect 8309 4505 8343 4539
rect 5733 4437 5767 4471
rect 6193 4437 6227 4471
rect 13277 4437 13311 4471
rect 15393 4437 15427 4471
rect 6561 4233 6595 4267
rect 8677 4233 8711 4267
rect 10517 4233 10551 4267
rect 12848 4165 12882 4199
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 7297 4097 7331 4131
rect 7564 4097 7598 4131
rect 9137 4097 9171 4131
rect 9404 4097 9438 4131
rect 13093 4097 13127 4131
rect 14861 4097 14895 4131
rect 15117 4097 15151 4131
rect 15577 4097 15611 4131
rect 13737 3961 13771 3995
rect 11713 3893 11747 3927
rect 15761 3893 15795 3927
rect 7481 3689 7515 3723
rect 9781 3689 9815 3723
rect 11253 3689 11287 3723
rect 6101 3553 6135 3587
rect 8953 3553 8987 3587
rect 10885 3553 10919 3587
rect 6357 3485 6391 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 11069 3485 11103 3519
rect 1593 2601 1627 2635
rect 1409 2397 1443 2431
rect 8953 2397 8987 2431
rect 16865 2397 16899 2431
rect 17049 2261 17083 2295
<< metal1 >>
rect 1104 47354 18860 47376
rect 1104 47302 3915 47354
rect 3967 47302 3979 47354
rect 4031 47302 4043 47354
rect 4095 47302 4107 47354
rect 4159 47302 4171 47354
rect 4223 47302 9846 47354
rect 9898 47302 9910 47354
rect 9962 47302 9974 47354
rect 10026 47302 10038 47354
rect 10090 47302 10102 47354
rect 10154 47302 15776 47354
rect 15828 47302 15840 47354
rect 15892 47302 15904 47354
rect 15956 47302 15968 47354
rect 16020 47302 16032 47354
rect 16084 47302 18860 47354
rect 1104 47280 18860 47302
rect 11054 47200 11060 47252
rect 11112 47240 11118 47252
rect 11517 47243 11575 47249
rect 11517 47240 11529 47243
rect 11112 47212 11529 47240
rect 11112 47200 11118 47212
rect 11517 47209 11529 47212
rect 11563 47209 11575 47243
rect 11517 47203 11575 47209
rect 18049 47243 18107 47249
rect 18049 47209 18061 47243
rect 18095 47240 18107 47243
rect 19334 47240 19340 47252
rect 18095 47212 19340 47240
rect 18095 47209 18107 47212
rect 18049 47203 18107 47209
rect 19334 47200 19340 47212
rect 19392 47200 19398 47252
rect 2774 47036 2780 47048
rect 2735 47008 2780 47036
rect 2774 46996 2780 47008
rect 2832 46996 2838 47048
rect 17862 47036 17868 47048
rect 17823 47008 17868 47036
rect 17862 46996 17868 47008
rect 17920 46996 17926 47048
rect 2961 46971 3019 46977
rect 2961 46937 2973 46971
rect 3007 46968 3019 46971
rect 3234 46968 3240 46980
rect 3007 46940 3240 46968
rect 3007 46937 3019 46940
rect 2961 46931 3019 46937
rect 3234 46928 3240 46940
rect 3292 46928 3298 46980
rect 1104 46810 18860 46832
rect 1104 46758 6880 46810
rect 6932 46758 6944 46810
rect 6996 46758 7008 46810
rect 7060 46758 7072 46810
rect 7124 46758 7136 46810
rect 7188 46758 12811 46810
rect 12863 46758 12875 46810
rect 12927 46758 12939 46810
rect 12991 46758 13003 46810
rect 13055 46758 13067 46810
rect 13119 46758 18860 46810
rect 1104 46736 18860 46758
rect 1104 46266 18860 46288
rect 1104 46214 3915 46266
rect 3967 46214 3979 46266
rect 4031 46214 4043 46266
rect 4095 46214 4107 46266
rect 4159 46214 4171 46266
rect 4223 46214 9846 46266
rect 9898 46214 9910 46266
rect 9962 46214 9974 46266
rect 10026 46214 10038 46266
rect 10090 46214 10102 46266
rect 10154 46214 15776 46266
rect 15828 46214 15840 46266
rect 15892 46214 15904 46266
rect 15956 46214 15968 46266
rect 16020 46214 16032 46266
rect 16084 46214 18860 46266
rect 1104 46192 18860 46214
rect 8846 45908 8852 45960
rect 8904 45948 8910 45960
rect 8941 45951 8999 45957
rect 8941 45948 8953 45951
rect 8904 45920 8953 45948
rect 8904 45908 8910 45920
rect 8941 45917 8953 45920
rect 8987 45917 8999 45951
rect 9122 45948 9128 45960
rect 9083 45920 9128 45948
rect 8941 45911 8999 45917
rect 9122 45908 9128 45920
rect 9180 45908 9186 45960
rect 9033 45815 9091 45821
rect 9033 45781 9045 45815
rect 9079 45812 9091 45815
rect 9214 45812 9220 45824
rect 9079 45784 9220 45812
rect 9079 45781 9091 45784
rect 9033 45775 9091 45781
rect 9214 45772 9220 45784
rect 9272 45772 9278 45824
rect 1104 45722 18860 45744
rect 1104 45670 6880 45722
rect 6932 45670 6944 45722
rect 6996 45670 7008 45722
rect 7060 45670 7072 45722
rect 7124 45670 7136 45722
rect 7188 45670 12811 45722
rect 12863 45670 12875 45722
rect 12927 45670 12939 45722
rect 12991 45670 13003 45722
rect 13055 45670 13067 45722
rect 13119 45670 18860 45722
rect 1104 45648 18860 45670
rect 8128 45580 8432 45608
rect 8128 45549 8156 45580
rect 6733 45543 6791 45549
rect 6733 45509 6745 45543
rect 6779 45540 6791 45543
rect 8113 45543 8171 45549
rect 6779 45512 7512 45540
rect 6779 45509 6791 45512
rect 6733 45503 6791 45509
rect 7484 45481 7512 45512
rect 8113 45509 8125 45543
rect 8159 45509 8171 45543
rect 8313 45543 8371 45549
rect 8313 45540 8325 45543
rect 8113 45503 8171 45509
rect 8312 45509 8325 45540
rect 8359 45509 8371 45543
rect 8312 45503 8371 45509
rect 7009 45475 7067 45481
rect 7009 45441 7021 45475
rect 7055 45441 7067 45475
rect 7009 45435 7067 45441
rect 7469 45475 7527 45481
rect 7469 45441 7481 45475
rect 7515 45441 7527 45475
rect 7469 45435 7527 45441
rect 7653 45475 7711 45481
rect 7653 45441 7665 45475
rect 7699 45472 7711 45475
rect 8312 45472 8340 45503
rect 7699 45444 8340 45472
rect 7699 45441 7711 45444
rect 7653 45435 7711 45441
rect 6178 45364 6184 45416
rect 6236 45404 6242 45416
rect 6733 45407 6791 45413
rect 6733 45404 6745 45407
rect 6236 45376 6745 45404
rect 6236 45364 6242 45376
rect 6733 45373 6745 45376
rect 6779 45373 6791 45407
rect 7024 45404 7052 45435
rect 8128 45416 8156 45444
rect 7926 45404 7932 45416
rect 7024 45376 7932 45404
rect 6733 45367 6791 45373
rect 7926 45364 7932 45376
rect 7984 45364 7990 45416
rect 8110 45364 8116 45416
rect 8168 45364 8174 45416
rect 8404 45404 8432 45580
rect 8846 45500 8852 45552
rect 8904 45540 8910 45552
rect 9953 45543 10011 45549
rect 8904 45512 9352 45540
rect 8904 45500 8910 45512
rect 9324 45481 9352 45512
rect 9953 45509 9965 45543
rect 9999 45540 10011 45543
rect 10318 45540 10324 45552
rect 9999 45512 10324 45540
rect 9999 45509 10011 45512
rect 9953 45503 10011 45509
rect 9125 45475 9183 45481
rect 9125 45441 9137 45475
rect 9171 45441 9183 45475
rect 9125 45435 9183 45441
rect 9309 45475 9367 45481
rect 9309 45441 9321 45475
rect 9355 45472 9367 45475
rect 9861 45475 9919 45481
rect 9861 45472 9873 45475
rect 9355 45444 9873 45472
rect 9355 45441 9367 45444
rect 9309 45435 9367 45441
rect 9861 45441 9873 45444
rect 9907 45441 9919 45475
rect 9861 45435 9919 45441
rect 9140 45404 9168 45435
rect 9401 45407 9459 45413
rect 8404 45376 9076 45404
rect 9140 45376 9352 45404
rect 8481 45339 8539 45345
rect 8481 45305 8493 45339
rect 8527 45336 8539 45339
rect 8846 45336 8852 45348
rect 8527 45308 8852 45336
rect 8527 45305 8539 45308
rect 8481 45299 8539 45305
rect 8846 45296 8852 45308
rect 8904 45296 8910 45348
rect 9048 45336 9076 45376
rect 9324 45336 9352 45376
rect 9401 45373 9413 45407
rect 9447 45404 9459 45407
rect 9968 45404 9996 45503
rect 10318 45500 10324 45512
rect 10376 45500 10382 45552
rect 10137 45475 10195 45481
rect 10137 45441 10149 45475
rect 10183 45472 10195 45475
rect 10410 45472 10416 45484
rect 10183 45444 10416 45472
rect 10183 45441 10195 45444
rect 10137 45435 10195 45441
rect 10410 45432 10416 45444
rect 10468 45432 10474 45484
rect 11514 45472 11520 45484
rect 11475 45444 11520 45472
rect 11514 45432 11520 45444
rect 11572 45432 11578 45484
rect 11701 45475 11759 45481
rect 11701 45441 11713 45475
rect 11747 45472 11759 45475
rect 12066 45472 12072 45484
rect 11747 45444 12072 45472
rect 11747 45441 11759 45444
rect 11701 45435 11759 45441
rect 12066 45432 12072 45444
rect 12124 45432 12130 45484
rect 9447 45376 9996 45404
rect 9447 45373 9459 45376
rect 9401 45367 9459 45373
rect 10137 45339 10195 45345
rect 10137 45336 10149 45339
rect 9048 45308 9260 45336
rect 9324 45308 10149 45336
rect 6914 45228 6920 45280
rect 6972 45268 6978 45280
rect 7466 45268 7472 45280
rect 6972 45240 7017 45268
rect 7427 45240 7472 45268
rect 6972 45228 6978 45240
rect 7466 45228 7472 45240
rect 7524 45228 7530 45280
rect 8297 45271 8355 45277
rect 8297 45237 8309 45271
rect 8343 45268 8355 45271
rect 8662 45268 8668 45280
rect 8343 45240 8668 45268
rect 8343 45237 8355 45240
rect 8297 45231 8355 45237
rect 8662 45228 8668 45240
rect 8720 45228 8726 45280
rect 8941 45271 8999 45277
rect 8941 45237 8953 45271
rect 8987 45268 8999 45271
rect 9030 45268 9036 45280
rect 8987 45240 9036 45268
rect 8987 45237 8999 45240
rect 8941 45231 8999 45237
rect 9030 45228 9036 45240
rect 9088 45228 9094 45280
rect 9232 45268 9260 45308
rect 10137 45305 10149 45308
rect 10183 45305 10195 45339
rect 10137 45299 10195 45305
rect 10226 45268 10232 45280
rect 9232 45240 10232 45268
rect 10226 45228 10232 45240
rect 10284 45228 10290 45280
rect 11517 45271 11575 45277
rect 11517 45237 11529 45271
rect 11563 45268 11575 45271
rect 13262 45268 13268 45280
rect 11563 45240 13268 45268
rect 11563 45237 11575 45240
rect 11517 45231 11575 45237
rect 13262 45228 13268 45240
rect 13320 45228 13326 45280
rect 1104 45178 18860 45200
rect 1104 45126 3915 45178
rect 3967 45126 3979 45178
rect 4031 45126 4043 45178
rect 4095 45126 4107 45178
rect 4159 45126 4171 45178
rect 4223 45126 9846 45178
rect 9898 45126 9910 45178
rect 9962 45126 9974 45178
rect 10026 45126 10038 45178
rect 10090 45126 10102 45178
rect 10154 45126 15776 45178
rect 15828 45126 15840 45178
rect 15892 45126 15904 45178
rect 15956 45126 15968 45178
rect 16020 45126 16032 45178
rect 16084 45126 18860 45178
rect 1104 45104 18860 45126
rect 6914 45024 6920 45076
rect 6972 45064 6978 45076
rect 7374 45064 7380 45076
rect 6972 45036 7380 45064
rect 6972 45024 6978 45036
rect 7374 45024 7380 45036
rect 7432 45024 7438 45076
rect 11517 44999 11575 45005
rect 11517 44965 11529 44999
rect 11563 44996 11575 44999
rect 17862 44996 17868 45008
rect 11563 44968 17868 44996
rect 11563 44965 11575 44968
rect 11517 44959 11575 44965
rect 17862 44956 17868 44968
rect 17920 44956 17926 45008
rect 5537 44863 5595 44869
rect 5537 44829 5549 44863
rect 5583 44860 5595 44863
rect 6362 44860 6368 44872
rect 5583 44832 6368 44860
rect 5583 44829 5595 44832
rect 5537 44823 5595 44829
rect 6362 44820 6368 44832
rect 6420 44820 6426 44872
rect 7558 44860 7564 44872
rect 7519 44832 7564 44860
rect 7558 44820 7564 44832
rect 7616 44820 7622 44872
rect 7653 44863 7711 44869
rect 7653 44829 7665 44863
rect 7699 44829 7711 44863
rect 7653 44823 7711 44829
rect 5810 44801 5816 44804
rect 5804 44755 5816 44801
rect 5868 44792 5874 44804
rect 7668 44792 7696 44823
rect 8018 44820 8024 44872
rect 8076 44860 8082 44872
rect 8205 44863 8263 44869
rect 8205 44860 8217 44863
rect 8076 44832 8217 44860
rect 8076 44820 8082 44832
rect 8205 44829 8217 44832
rect 8251 44829 8263 44863
rect 8205 44823 8263 44829
rect 5868 44764 5904 44792
rect 6932 44764 7696 44792
rect 8220 44792 8248 44823
rect 8294 44820 8300 44872
rect 8352 44860 8358 44872
rect 8389 44863 8447 44869
rect 8389 44860 8401 44863
rect 8352 44832 8401 44860
rect 8352 44820 8358 44832
rect 8389 44829 8401 44832
rect 8435 44829 8447 44863
rect 8938 44860 8944 44872
rect 8899 44832 8944 44860
rect 8389 44823 8447 44829
rect 8938 44820 8944 44832
rect 8996 44820 9002 44872
rect 9030 44820 9036 44872
rect 9088 44860 9094 44872
rect 9197 44863 9255 44869
rect 9197 44860 9209 44863
rect 9088 44832 9209 44860
rect 9088 44820 9094 44832
rect 9197 44829 9209 44832
rect 9243 44829 9255 44863
rect 10870 44860 10876 44872
rect 10831 44832 10876 44860
rect 9197 44823 9255 44829
rect 10870 44820 10876 44832
rect 10928 44820 10934 44872
rect 11149 44863 11207 44869
rect 11149 44829 11161 44863
rect 11195 44829 11207 44863
rect 11422 44860 11428 44872
rect 11383 44832 11428 44860
rect 11149 44823 11207 44829
rect 10410 44792 10416 44804
rect 8220 44764 10416 44792
rect 5810 44752 5816 44755
rect 5868 44752 5874 44764
rect 6546 44684 6552 44736
rect 6604 44724 6610 44736
rect 6932 44733 6960 44764
rect 10410 44752 10416 44764
rect 10468 44752 10474 44804
rect 11164 44792 11192 44823
rect 11422 44820 11428 44832
rect 11480 44820 11486 44872
rect 11606 44860 11612 44872
rect 11567 44832 11612 44860
rect 11606 44820 11612 44832
rect 11664 44820 11670 44872
rect 12066 44860 12072 44872
rect 12027 44832 12072 44860
rect 12066 44820 12072 44832
rect 12124 44820 12130 44872
rect 11330 44792 11336 44804
rect 11164 44764 11336 44792
rect 11330 44752 11336 44764
rect 11388 44792 11394 44804
rect 12161 44795 12219 44801
rect 12161 44792 12173 44795
rect 11388 44764 12173 44792
rect 11388 44752 11394 44764
rect 12161 44761 12173 44764
rect 12207 44761 12219 44795
rect 12161 44755 12219 44761
rect 6917 44727 6975 44733
rect 6917 44724 6929 44727
rect 6604 44696 6929 44724
rect 6604 44684 6610 44696
rect 6917 44693 6929 44696
rect 6963 44693 6975 44727
rect 6917 44687 6975 44693
rect 8297 44727 8355 44733
rect 8297 44693 8309 44727
rect 8343 44724 8355 44727
rect 8386 44724 8392 44736
rect 8343 44696 8392 44724
rect 8343 44693 8355 44696
rect 8297 44687 8355 44693
rect 8386 44684 8392 44696
rect 8444 44684 8450 44736
rect 10318 44724 10324 44736
rect 10231 44696 10324 44724
rect 10318 44684 10324 44696
rect 10376 44724 10382 44736
rect 10870 44724 10876 44736
rect 10376 44696 10876 44724
rect 10376 44684 10382 44696
rect 10870 44684 10876 44696
rect 10928 44684 10934 44736
rect 1104 44634 18860 44656
rect 1104 44582 6880 44634
rect 6932 44582 6944 44634
rect 6996 44582 7008 44634
rect 7060 44582 7072 44634
rect 7124 44582 7136 44634
rect 7188 44582 12811 44634
rect 12863 44582 12875 44634
rect 12927 44582 12939 44634
rect 12991 44582 13003 44634
rect 13055 44582 13067 44634
rect 13119 44582 18860 44634
rect 1104 44560 18860 44582
rect 5721 44523 5779 44529
rect 5721 44489 5733 44523
rect 5767 44520 5779 44523
rect 5810 44520 5816 44532
rect 5767 44492 5816 44520
rect 5767 44489 5779 44492
rect 5721 44483 5779 44489
rect 5810 44480 5816 44492
rect 5868 44480 5874 44532
rect 6365 44523 6423 44529
rect 6365 44489 6377 44523
rect 6411 44520 6423 44523
rect 7926 44520 7932 44532
rect 6411 44492 7932 44520
rect 6411 44489 6423 44492
rect 6365 44483 6423 44489
rect 7926 44480 7932 44492
rect 7984 44480 7990 44532
rect 11517 44523 11575 44529
rect 11517 44489 11529 44523
rect 11563 44520 11575 44523
rect 12066 44520 12072 44532
rect 11563 44492 12072 44520
rect 11563 44489 11575 44492
rect 11517 44483 11575 44489
rect 12066 44480 12072 44492
rect 12124 44480 12130 44532
rect 7374 44452 7380 44464
rect 5644 44424 7380 44452
rect 1854 44384 1860 44396
rect 1815 44356 1860 44384
rect 1854 44344 1860 44356
rect 1912 44344 1918 44396
rect 5644 44393 5672 44424
rect 7374 44412 7380 44424
rect 7432 44412 7438 44464
rect 7466 44412 7472 44464
rect 7524 44461 7530 44464
rect 7524 44452 7536 44461
rect 7524 44424 7569 44452
rect 10980 44424 12940 44452
rect 7524 44415 7536 44424
rect 7524 44412 7530 44415
rect 5629 44387 5687 44393
rect 5629 44353 5641 44387
rect 5675 44353 5687 44387
rect 5810 44384 5816 44396
rect 5771 44356 5816 44384
rect 5629 44347 5687 44353
rect 5810 44344 5816 44356
rect 5868 44344 5874 44396
rect 7834 44384 7840 44396
rect 5920 44356 7840 44384
rect 2133 44319 2191 44325
rect 2133 44285 2145 44319
rect 2179 44316 2191 44319
rect 5920 44316 5948 44356
rect 7834 44344 7840 44356
rect 7892 44344 7898 44396
rect 8386 44384 8392 44396
rect 8347 44356 8392 44384
rect 8386 44344 8392 44356
rect 8444 44344 8450 44396
rect 8662 44384 8668 44396
rect 8623 44356 8668 44384
rect 8662 44344 8668 44356
rect 8720 44344 8726 44396
rect 10318 44344 10324 44396
rect 10376 44384 10382 44396
rect 10980 44393 11008 44424
rect 10698 44387 10756 44393
rect 10698 44384 10710 44387
rect 10376 44356 10710 44384
rect 10376 44344 10382 44356
rect 10698 44353 10710 44356
rect 10744 44353 10756 44387
rect 10698 44347 10756 44353
rect 10965 44387 11023 44393
rect 10965 44353 10977 44387
rect 11011 44353 11023 44387
rect 10965 44347 11023 44353
rect 12641 44387 12699 44393
rect 12641 44353 12653 44387
rect 12687 44384 12699 44387
rect 12802 44384 12808 44396
rect 12687 44356 12808 44384
rect 12687 44353 12699 44356
rect 12641 44347 12699 44353
rect 12802 44344 12808 44356
rect 12860 44344 12866 44396
rect 12912 44393 12940 44424
rect 12897 44387 12955 44393
rect 12897 44353 12909 44387
rect 12943 44384 12955 44387
rect 13814 44384 13820 44396
rect 12943 44356 13820 44384
rect 12943 44353 12955 44356
rect 12897 44347 12955 44353
rect 13814 44344 13820 44356
rect 13872 44344 13878 44396
rect 7742 44316 7748 44328
rect 2179 44288 5948 44316
rect 7703 44288 7748 44316
rect 2179 44285 2191 44288
rect 2133 44279 2191 44285
rect 7742 44276 7748 44288
rect 7800 44276 7806 44328
rect 8110 44208 8116 44260
rect 8168 44248 8174 44260
rect 8573 44251 8631 44257
rect 8573 44248 8585 44251
rect 8168 44220 8585 44248
rect 8168 44208 8174 44220
rect 8573 44217 8585 44220
rect 8619 44217 8631 44251
rect 8573 44211 8631 44217
rect 7466 44140 7472 44192
rect 7524 44180 7530 44192
rect 8205 44183 8263 44189
rect 8205 44180 8217 44183
rect 7524 44152 8217 44180
rect 7524 44140 7530 44152
rect 8205 44149 8217 44152
rect 8251 44149 8263 44183
rect 8205 44143 8263 44149
rect 9585 44183 9643 44189
rect 9585 44149 9597 44183
rect 9631 44180 9643 44183
rect 9766 44180 9772 44192
rect 9631 44152 9772 44180
rect 9631 44149 9643 44152
rect 9585 44143 9643 44149
rect 9766 44140 9772 44152
rect 9824 44140 9830 44192
rect 1104 44090 18860 44112
rect 1104 44038 3915 44090
rect 3967 44038 3979 44090
rect 4031 44038 4043 44090
rect 4095 44038 4107 44090
rect 4159 44038 4171 44090
rect 4223 44038 9846 44090
rect 9898 44038 9910 44090
rect 9962 44038 9974 44090
rect 10026 44038 10038 44090
rect 10090 44038 10102 44090
rect 10154 44038 15776 44090
rect 15828 44038 15840 44090
rect 15892 44038 15904 44090
rect 15956 44038 15968 44090
rect 16020 44038 16032 44090
rect 16084 44038 18860 44090
rect 1104 44016 18860 44038
rect 5810 43936 5816 43988
rect 5868 43976 5874 43988
rect 6273 43979 6331 43985
rect 6273 43976 6285 43979
rect 5868 43948 6285 43976
rect 5868 43936 5874 43948
rect 6273 43945 6285 43948
rect 6319 43945 6331 43979
rect 7558 43976 7564 43988
rect 6273 43939 6331 43945
rect 6886 43948 7564 43976
rect 6365 43911 6423 43917
rect 6365 43877 6377 43911
rect 6411 43908 6423 43911
rect 6454 43908 6460 43920
rect 6411 43880 6460 43908
rect 6411 43877 6423 43880
rect 6365 43871 6423 43877
rect 6454 43868 6460 43880
rect 6512 43908 6518 43920
rect 6886 43908 6914 43948
rect 7558 43936 7564 43948
rect 7616 43936 7622 43988
rect 8297 43979 8355 43985
rect 8297 43945 8309 43979
rect 8343 43976 8355 43979
rect 8662 43976 8668 43988
rect 8343 43948 8668 43976
rect 8343 43945 8355 43948
rect 8297 43939 8355 43945
rect 8662 43936 8668 43948
rect 8720 43936 8726 43988
rect 10226 43936 10232 43988
rect 10284 43976 10290 43988
rect 10321 43979 10379 43985
rect 10321 43976 10333 43979
rect 10284 43948 10333 43976
rect 10284 43936 10290 43948
rect 10321 43945 10333 43948
rect 10367 43945 10379 43979
rect 10321 43939 10379 43945
rect 11422 43936 11428 43988
rect 11480 43976 11486 43988
rect 11517 43979 11575 43985
rect 11517 43976 11529 43979
rect 11480 43948 11529 43976
rect 11480 43936 11486 43948
rect 11517 43945 11529 43948
rect 11563 43945 11575 43979
rect 11517 43939 11575 43945
rect 12802 43936 12808 43988
rect 12860 43976 12866 43988
rect 13357 43979 13415 43985
rect 13357 43976 13369 43979
rect 12860 43948 13369 43976
rect 12860 43936 12866 43948
rect 13357 43945 13369 43948
rect 13403 43945 13415 43979
rect 13357 43939 13415 43945
rect 6512 43880 6914 43908
rect 6512 43868 6518 43880
rect 11606 43868 11612 43920
rect 11664 43908 11670 43920
rect 13262 43908 13268 43920
rect 11664 43880 12388 43908
rect 13223 43880 13268 43908
rect 11664 43868 11670 43880
rect 6178 43840 6184 43852
rect 6139 43812 6184 43840
rect 6178 43800 6184 43812
rect 6236 43800 6242 43852
rect 6917 43843 6975 43849
rect 6917 43840 6929 43843
rect 6380 43812 6929 43840
rect 6380 43784 6408 43812
rect 6917 43809 6929 43812
rect 6963 43809 6975 43843
rect 6917 43803 6975 43809
rect 6362 43732 6368 43784
rect 6420 43732 6426 43784
rect 6457 43775 6515 43781
rect 6457 43741 6469 43775
rect 6503 43772 6515 43775
rect 6546 43772 6552 43784
rect 6503 43744 6552 43772
rect 6503 43741 6515 43744
rect 6457 43735 6515 43741
rect 6546 43732 6552 43744
rect 6604 43732 6610 43784
rect 6932 43704 6960 43803
rect 10870 43800 10876 43852
rect 10928 43840 10934 43852
rect 11149 43843 11207 43849
rect 11149 43840 11161 43843
rect 10928 43812 11161 43840
rect 10928 43800 10934 43812
rect 11149 43809 11161 43812
rect 11195 43809 11207 43843
rect 12250 43840 12256 43852
rect 12211 43812 12256 43840
rect 11149 43803 11207 43809
rect 12250 43800 12256 43812
rect 12308 43800 12314 43852
rect 12360 43840 12388 43880
rect 13262 43868 13268 43880
rect 13320 43868 13326 43920
rect 13357 43843 13415 43849
rect 13357 43840 13369 43843
rect 12360 43812 13369 43840
rect 13357 43809 13369 43812
rect 13403 43809 13415 43843
rect 13357 43803 13415 43809
rect 7184 43775 7242 43781
rect 7184 43741 7196 43775
rect 7230 43774 7242 43775
rect 7230 43772 7328 43774
rect 7466 43772 7472 43784
rect 7230 43746 7472 43772
rect 7230 43741 7242 43746
rect 7300 43744 7472 43746
rect 7184 43735 7242 43741
rect 7466 43732 7472 43744
rect 7524 43732 7530 43784
rect 7742 43732 7748 43784
rect 7800 43772 7806 43784
rect 8938 43772 8944 43784
rect 7800 43744 8944 43772
rect 7800 43732 7806 43744
rect 8938 43732 8944 43744
rect 8996 43732 9002 43784
rect 9214 43781 9220 43784
rect 9208 43735 9220 43781
rect 9272 43772 9278 43784
rect 10778 43772 10784 43784
rect 9272 43744 9308 43772
rect 10739 43744 10784 43772
rect 9214 43732 9220 43735
rect 9272 43732 9278 43744
rect 10778 43732 10784 43744
rect 10836 43732 10842 43784
rect 10965 43775 11023 43781
rect 10965 43741 10977 43775
rect 11011 43741 11023 43775
rect 10965 43735 11023 43741
rect 11057 43775 11115 43781
rect 11057 43741 11069 43775
rect 11103 43741 11115 43775
rect 11330 43772 11336 43784
rect 11291 43744 11336 43772
rect 11057 43735 11115 43741
rect 7760 43704 7788 43732
rect 6932 43676 7788 43704
rect 10226 43664 10232 43716
rect 10284 43704 10290 43716
rect 10980 43704 11008 43735
rect 10284 43676 11008 43704
rect 10284 43664 10290 43676
rect 10962 43596 10968 43648
rect 11020 43636 11026 43648
rect 11072 43636 11100 43735
rect 11330 43732 11336 43744
rect 11388 43772 11394 43784
rect 12345 43775 12403 43781
rect 12345 43772 12357 43775
rect 11388 43744 12357 43772
rect 11388 43732 11394 43744
rect 12345 43741 12357 43744
rect 12391 43741 12403 43775
rect 12345 43735 12403 43741
rect 12434 43664 12440 43716
rect 12492 43704 12498 43716
rect 12989 43707 13047 43713
rect 12989 43704 13001 43707
rect 12492 43676 13001 43704
rect 12492 43664 12498 43676
rect 12989 43673 13001 43676
rect 13035 43673 13047 43707
rect 12989 43667 13047 43673
rect 11974 43636 11980 43648
rect 11020 43608 11100 43636
rect 11935 43608 11980 43636
rect 11020 43596 11026 43608
rect 11974 43596 11980 43608
rect 12032 43596 12038 43648
rect 12526 43596 12532 43648
rect 12584 43636 12590 43648
rect 13081 43639 13139 43645
rect 13081 43636 13093 43639
rect 12584 43608 13093 43636
rect 12584 43596 12590 43608
rect 13081 43605 13093 43608
rect 13127 43636 13139 43639
rect 13262 43636 13268 43648
rect 13127 43608 13268 43636
rect 13127 43605 13139 43608
rect 13081 43599 13139 43605
rect 13262 43596 13268 43608
rect 13320 43596 13326 43648
rect 1104 43546 18860 43568
rect 1104 43494 6880 43546
rect 6932 43494 6944 43546
rect 6996 43494 7008 43546
rect 7060 43494 7072 43546
rect 7124 43494 7136 43546
rect 7188 43494 12811 43546
rect 12863 43494 12875 43546
rect 12927 43494 12939 43546
rect 12991 43494 13003 43546
rect 13055 43494 13067 43546
rect 13119 43494 18860 43546
rect 1104 43472 18860 43494
rect 6454 43392 6460 43444
rect 6512 43432 6518 43444
rect 7209 43435 7267 43441
rect 7209 43432 7221 43435
rect 6512 43404 7221 43432
rect 6512 43392 6518 43404
rect 7209 43401 7221 43404
rect 7255 43401 7267 43435
rect 7209 43395 7267 43401
rect 9861 43435 9919 43441
rect 9861 43401 9873 43435
rect 9907 43432 9919 43435
rect 10778 43432 10784 43444
rect 9907 43404 10784 43432
rect 9907 43401 9919 43404
rect 9861 43395 9919 43401
rect 10778 43392 10784 43404
rect 10836 43392 10842 43444
rect 12434 43432 12440 43444
rect 12395 43404 12440 43432
rect 12434 43392 12440 43404
rect 12492 43392 12498 43444
rect 7009 43367 7067 43373
rect 7009 43333 7021 43367
rect 7055 43364 7067 43367
rect 7926 43364 7932 43376
rect 7055 43336 7932 43364
rect 7055 43333 7067 43336
rect 7009 43327 7067 43333
rect 7926 43324 7932 43336
rect 7984 43364 7990 43376
rect 8570 43364 8576 43376
rect 7984 43336 8576 43364
rect 7984 43324 7990 43336
rect 8570 43324 8576 43336
rect 8628 43324 8634 43376
rect 9493 43367 9551 43373
rect 9493 43364 9505 43367
rect 8680 43336 9505 43364
rect 8680 43308 8708 43336
rect 9493 43333 9505 43336
rect 9539 43333 9551 43367
rect 9493 43327 9551 43333
rect 9585 43367 9643 43373
rect 9585 43333 9597 43367
rect 9631 43364 9643 43367
rect 10318 43364 10324 43376
rect 9631 43336 10180 43364
rect 10279 43336 10324 43364
rect 9631 43333 9643 43336
rect 9585 43327 9643 43333
rect 8110 43296 8116 43308
rect 7392 43268 8116 43296
rect 7392 43169 7420 43268
rect 8110 43256 8116 43268
rect 8168 43256 8174 43308
rect 8297 43299 8355 43305
rect 8297 43265 8309 43299
rect 8343 43296 8355 43299
rect 8662 43296 8668 43308
rect 8343 43268 8668 43296
rect 8343 43265 8355 43268
rect 8297 43259 8355 43265
rect 8662 43256 8668 43268
rect 8720 43256 8726 43308
rect 9214 43296 9220 43308
rect 9175 43268 9220 43296
rect 9214 43256 9220 43268
rect 9272 43256 9278 43308
rect 9365 43299 9423 43305
rect 9365 43265 9377 43299
rect 9411 43296 9423 43299
rect 9674 43296 9680 43308
rect 9732 43305 9738 43308
rect 9411 43265 9444 43296
rect 9592 43268 9680 43296
rect 9365 43259 9444 43265
rect 9416 43228 9444 43259
rect 9674 43256 9680 43268
rect 9732 43296 9740 43305
rect 10152 43296 10180 43336
rect 10318 43324 10324 43336
rect 10376 43324 10382 43376
rect 10962 43364 10968 43376
rect 10520 43336 10968 43364
rect 10520 43296 10548 43336
rect 10962 43324 10968 43336
rect 11020 43324 11026 43376
rect 9732 43268 9812 43296
rect 10152 43268 10548 43296
rect 10689 43299 10747 43305
rect 9732 43259 9740 43268
rect 9732 43256 9738 43259
rect 9784 43228 9812 43268
rect 10689 43265 10701 43299
rect 10735 43265 10747 43299
rect 10689 43259 10747 43265
rect 10226 43228 10232 43240
rect 9416 43200 9628 43228
rect 9784 43200 10232 43228
rect 9600 43172 9628 43200
rect 10226 43188 10232 43200
rect 10284 43188 10290 43240
rect 10413 43231 10471 43237
rect 10413 43197 10425 43231
rect 10459 43228 10471 43231
rect 10704 43228 10732 43259
rect 10778 43256 10784 43308
rect 10836 43296 10842 43308
rect 10836 43268 10881 43296
rect 10836 43256 10842 43268
rect 11882 43256 11888 43308
rect 11940 43296 11946 43308
rect 12069 43299 12127 43305
rect 12069 43296 12081 43299
rect 11940 43268 12081 43296
rect 11940 43256 11946 43268
rect 12069 43265 12081 43268
rect 12115 43265 12127 43299
rect 12069 43259 12127 43265
rect 11974 43228 11980 43240
rect 10459 43200 10640 43228
rect 10704 43200 10824 43228
rect 11935 43200 11980 43228
rect 10459 43197 10471 43200
rect 10413 43191 10471 43197
rect 7377 43163 7435 43169
rect 7377 43129 7389 43163
rect 7423 43129 7435 43163
rect 7377 43123 7435 43129
rect 9582 43120 9588 43172
rect 9640 43120 9646 43172
rect 6546 43052 6552 43104
rect 6604 43092 6610 43104
rect 7193 43095 7251 43101
rect 7193 43092 7205 43095
rect 6604 43064 7205 43092
rect 6604 43052 6610 43064
rect 7193 43061 7205 43064
rect 7239 43092 7251 43095
rect 7742 43092 7748 43104
rect 7239 43064 7748 43092
rect 7239 43061 7251 43064
rect 7193 43055 7251 43061
rect 7742 43052 7748 43064
rect 7800 43052 7806 43104
rect 7929 43095 7987 43101
rect 7929 43061 7941 43095
rect 7975 43092 7987 43095
rect 8294 43092 8300 43104
rect 7975 43064 8300 43092
rect 7975 43061 7987 43064
rect 7929 43055 7987 43061
rect 8294 43052 8300 43064
rect 8352 43052 8358 43104
rect 10502 43092 10508 43104
rect 10463 43064 10508 43092
rect 10502 43052 10508 43064
rect 10560 43052 10566 43104
rect 10612 43092 10640 43200
rect 10796 43160 10824 43200
rect 11974 43188 11980 43200
rect 12032 43188 12038 43240
rect 12526 43160 12532 43172
rect 10796 43132 12532 43160
rect 12526 43120 12532 43132
rect 12584 43120 12590 43172
rect 10870 43092 10876 43104
rect 10612 43064 10876 43092
rect 10870 43052 10876 43064
rect 10928 43092 10934 43104
rect 11606 43092 11612 43104
rect 10928 43064 11612 43092
rect 10928 43052 10934 43064
rect 11606 43052 11612 43064
rect 11664 43052 11670 43104
rect 1104 43002 18860 43024
rect 1104 42950 3915 43002
rect 3967 42950 3979 43002
rect 4031 42950 4043 43002
rect 4095 42950 4107 43002
rect 4159 42950 4171 43002
rect 4223 42950 9846 43002
rect 9898 42950 9910 43002
rect 9962 42950 9974 43002
rect 10026 42950 10038 43002
rect 10090 42950 10102 43002
rect 10154 42950 15776 43002
rect 15828 42950 15840 43002
rect 15892 42950 15904 43002
rect 15956 42950 15968 43002
rect 16020 42950 16032 43002
rect 16084 42950 18860 43002
rect 1104 42928 18860 42950
rect 8294 42848 8300 42900
rect 8352 42888 8358 42900
rect 9125 42891 9183 42897
rect 9125 42888 9137 42891
rect 8352 42860 9137 42888
rect 8352 42848 8358 42860
rect 9125 42857 9137 42860
rect 9171 42857 9183 42891
rect 9125 42851 9183 42857
rect 6178 42780 6184 42832
rect 6236 42820 6242 42832
rect 6236 42792 8984 42820
rect 6236 42780 6242 42792
rect 8956 42761 8984 42792
rect 8941 42755 8999 42761
rect 8941 42721 8953 42755
rect 8987 42752 8999 42755
rect 9030 42752 9036 42764
rect 8987 42724 9036 42752
rect 8987 42721 8999 42724
rect 8941 42715 8999 42721
rect 9030 42712 9036 42724
rect 9088 42712 9094 42764
rect 10962 42752 10968 42764
rect 10923 42724 10968 42752
rect 10962 42712 10968 42724
rect 11020 42712 11026 42764
rect 9217 42687 9275 42693
rect 9217 42653 9229 42687
rect 9263 42684 9275 42687
rect 9674 42684 9680 42696
rect 9263 42656 9680 42684
rect 9263 42653 9275 42656
rect 9217 42647 9275 42653
rect 9674 42644 9680 42656
rect 9732 42644 9738 42696
rect 9766 42644 9772 42696
rect 9824 42684 9830 42696
rect 9861 42687 9919 42693
rect 9861 42684 9873 42687
rect 9824 42656 9873 42684
rect 9824 42644 9830 42656
rect 9861 42653 9873 42656
rect 9907 42653 9919 42687
rect 9861 42647 9919 42653
rect 11057 42687 11115 42693
rect 11057 42653 11069 42687
rect 11103 42684 11115 42687
rect 12434 42684 12440 42696
rect 11103 42656 12440 42684
rect 11103 42653 11115 42656
rect 11057 42647 11115 42653
rect 12434 42644 12440 42656
rect 12492 42644 12498 42696
rect 8941 42551 8999 42557
rect 8941 42517 8953 42551
rect 8987 42548 8999 42551
rect 9122 42548 9128 42560
rect 8987 42520 9128 42548
rect 8987 42517 8999 42520
rect 8941 42511 8999 42517
rect 9122 42508 9128 42520
rect 9180 42508 9186 42560
rect 9582 42508 9588 42560
rect 9640 42548 9646 42560
rect 9769 42551 9827 42557
rect 9769 42548 9781 42551
rect 9640 42520 9781 42548
rect 9640 42508 9646 42520
rect 9769 42517 9781 42520
rect 9815 42517 9827 42551
rect 9769 42511 9827 42517
rect 1104 42458 18860 42480
rect 1104 42406 6880 42458
rect 6932 42406 6944 42458
rect 6996 42406 7008 42458
rect 7060 42406 7072 42458
rect 7124 42406 7136 42458
rect 7188 42406 12811 42458
rect 12863 42406 12875 42458
rect 12927 42406 12939 42458
rect 12991 42406 13003 42458
rect 13055 42406 13067 42458
rect 13119 42406 18860 42458
rect 1104 42384 18860 42406
rect 9125 42347 9183 42353
rect 9125 42313 9137 42347
rect 9171 42344 9183 42347
rect 9214 42344 9220 42356
rect 9171 42316 9220 42344
rect 9171 42313 9183 42316
rect 9125 42307 9183 42313
rect 9214 42304 9220 42316
rect 9272 42304 9278 42356
rect 10321 42347 10379 42353
rect 10321 42313 10333 42347
rect 10367 42344 10379 42347
rect 10502 42344 10508 42356
rect 10367 42316 10508 42344
rect 10367 42313 10379 42316
rect 10321 42307 10379 42313
rect 10502 42304 10508 42316
rect 10560 42304 10566 42356
rect 8662 42236 8668 42288
rect 8720 42276 8726 42288
rect 8720 42248 8800 42276
rect 8720 42236 8726 42248
rect 7561 42211 7619 42217
rect 7561 42177 7573 42211
rect 7607 42208 7619 42211
rect 7650 42208 7656 42220
rect 7607 42180 7656 42208
rect 7607 42177 7619 42180
rect 7561 42171 7619 42177
rect 7650 42168 7656 42180
rect 7708 42208 7714 42220
rect 7834 42208 7840 42220
rect 7708 42180 7840 42208
rect 7708 42168 7714 42180
rect 7834 42168 7840 42180
rect 7892 42168 7898 42220
rect 8386 42208 8392 42220
rect 8347 42180 8392 42208
rect 8386 42168 8392 42180
rect 8444 42168 8450 42220
rect 8570 42208 8576 42220
rect 8531 42180 8576 42208
rect 8570 42168 8576 42180
rect 8628 42168 8634 42220
rect 8772 42217 8800 42248
rect 8757 42211 8815 42217
rect 8757 42177 8769 42211
rect 8803 42177 8815 42211
rect 8757 42171 8815 42177
rect 8941 42211 8999 42217
rect 8941 42177 8953 42211
rect 8987 42208 8999 42211
rect 9582 42208 9588 42220
rect 8987 42180 9588 42208
rect 8987 42177 8999 42180
rect 8941 42171 8999 42177
rect 9582 42168 9588 42180
rect 9640 42168 9646 42220
rect 9766 42168 9772 42220
rect 9824 42208 9830 42220
rect 10229 42211 10287 42217
rect 10229 42208 10241 42211
rect 9824 42180 10241 42208
rect 9824 42168 9830 42180
rect 10229 42177 10241 42180
rect 10275 42177 10287 42211
rect 10229 42171 10287 42177
rect 10413 42211 10471 42217
rect 10413 42177 10425 42211
rect 10459 42208 10471 42211
rect 10870 42208 10876 42220
rect 10459 42180 10876 42208
rect 10459 42177 10471 42180
rect 10413 42171 10471 42177
rect 10870 42168 10876 42180
rect 10928 42208 10934 42220
rect 11514 42208 11520 42220
rect 10928 42180 11520 42208
rect 10928 42168 10934 42180
rect 11514 42168 11520 42180
rect 11572 42168 11578 42220
rect 8478 42100 8484 42152
rect 8536 42140 8542 42152
rect 8665 42143 8723 42149
rect 8665 42140 8677 42143
rect 8536 42112 8677 42140
rect 8536 42100 8542 42112
rect 8665 42109 8677 42112
rect 8711 42109 8723 42143
rect 8665 42103 8723 42109
rect 7837 42007 7895 42013
rect 7837 41973 7849 42007
rect 7883 42004 7895 42007
rect 7926 42004 7932 42016
rect 7883 41976 7932 42004
rect 7883 41973 7895 41976
rect 7837 41967 7895 41973
rect 7926 41964 7932 41976
rect 7984 41964 7990 42016
rect 1104 41914 18860 41936
rect 1104 41862 3915 41914
rect 3967 41862 3979 41914
rect 4031 41862 4043 41914
rect 4095 41862 4107 41914
rect 4159 41862 4171 41914
rect 4223 41862 9846 41914
rect 9898 41862 9910 41914
rect 9962 41862 9974 41914
rect 10026 41862 10038 41914
rect 10090 41862 10102 41914
rect 10154 41862 15776 41914
rect 15828 41862 15840 41914
rect 15892 41862 15904 41914
rect 15956 41862 15968 41914
rect 16020 41862 16032 41914
rect 16084 41862 18860 41914
rect 1104 41840 18860 41862
rect 1104 41370 18860 41392
rect 1104 41318 6880 41370
rect 6932 41318 6944 41370
rect 6996 41318 7008 41370
rect 7060 41318 7072 41370
rect 7124 41318 7136 41370
rect 7188 41318 12811 41370
rect 12863 41318 12875 41370
rect 12927 41318 12939 41370
rect 12991 41318 13003 41370
rect 13055 41318 13067 41370
rect 13119 41318 18860 41370
rect 1104 41296 18860 41318
rect 8386 41216 8392 41268
rect 8444 41256 8450 41268
rect 8665 41259 8723 41265
rect 8665 41256 8677 41259
rect 8444 41228 8677 41256
rect 8444 41216 8450 41228
rect 8665 41225 8677 41228
rect 8711 41225 8723 41259
rect 8665 41219 8723 41225
rect 8294 41188 8300 41200
rect 8255 41160 8300 41188
rect 8294 41148 8300 41160
rect 8352 41148 8358 41200
rect 8110 41120 8116 41132
rect 8071 41092 8116 41120
rect 8110 41080 8116 41092
rect 8168 41080 8174 41132
rect 8386 41120 8392 41132
rect 8347 41092 8392 41120
rect 8386 41080 8392 41092
rect 8444 41080 8450 41132
rect 8481 41123 8539 41129
rect 8481 41089 8493 41123
rect 8527 41120 8539 41123
rect 8570 41120 8576 41132
rect 8527 41092 8576 41120
rect 8527 41089 8539 41092
rect 8481 41083 8539 41089
rect 8570 41080 8576 41092
rect 8628 41080 8634 41132
rect 14645 41123 14703 41129
rect 14645 41089 14657 41123
rect 14691 41089 14703 41123
rect 14645 41083 14703 41089
rect 14829 41123 14887 41129
rect 14829 41089 14841 41123
rect 14875 41120 14887 41123
rect 15289 41123 15347 41129
rect 15289 41120 15301 41123
rect 14875 41092 15301 41120
rect 14875 41089 14887 41092
rect 14829 41083 14887 41089
rect 15289 41089 15301 41092
rect 15335 41089 15347 41123
rect 15289 41083 15347 41089
rect 15933 41123 15991 41129
rect 15933 41089 15945 41123
rect 15979 41120 15991 41123
rect 16666 41120 16672 41132
rect 15979 41092 16672 41120
rect 15979 41089 15991 41092
rect 15933 41083 15991 41089
rect 14458 41052 14464 41064
rect 14419 41024 14464 41052
rect 14458 41012 14464 41024
rect 14516 41012 14522 41064
rect 14660 41052 14688 41083
rect 16666 41080 16672 41092
rect 16724 41080 16730 41132
rect 18138 41120 18144 41132
rect 18099 41092 18144 41120
rect 18138 41080 18144 41092
rect 18196 41080 18202 41132
rect 15378 41052 15384 41064
rect 14660 41024 15384 41052
rect 15378 41012 15384 41024
rect 15436 41012 15442 41064
rect 15470 40916 15476 40928
rect 15431 40888 15476 40916
rect 15470 40876 15476 40888
rect 15528 40876 15534 40928
rect 16114 40916 16120 40928
rect 16075 40888 16120 40916
rect 16114 40876 16120 40888
rect 16172 40876 16178 40928
rect 17954 40916 17960 40928
rect 17915 40888 17960 40916
rect 17954 40876 17960 40888
rect 18012 40876 18018 40928
rect 1104 40826 18860 40848
rect 1104 40774 3915 40826
rect 3967 40774 3979 40826
rect 4031 40774 4043 40826
rect 4095 40774 4107 40826
rect 4159 40774 4171 40826
rect 4223 40774 9846 40826
rect 9898 40774 9910 40826
rect 9962 40774 9974 40826
rect 10026 40774 10038 40826
rect 10090 40774 10102 40826
rect 10154 40774 15776 40826
rect 15828 40774 15840 40826
rect 15892 40774 15904 40826
rect 15956 40774 15968 40826
rect 16020 40774 16032 40826
rect 16084 40774 18860 40826
rect 1104 40752 18860 40774
rect 6638 40672 6644 40724
rect 6696 40712 6702 40724
rect 6825 40715 6883 40721
rect 6825 40712 6837 40715
rect 6696 40684 6837 40712
rect 6696 40672 6702 40684
rect 6825 40681 6837 40684
rect 6871 40681 6883 40715
rect 8294 40712 8300 40724
rect 8255 40684 8300 40712
rect 6825 40675 6883 40681
rect 8294 40672 8300 40684
rect 8352 40672 8358 40724
rect 8386 40672 8392 40724
rect 8444 40712 8450 40724
rect 9125 40715 9183 40721
rect 9125 40712 9137 40715
rect 8444 40684 9137 40712
rect 8444 40672 8450 40684
rect 9125 40681 9137 40684
rect 9171 40681 9183 40715
rect 9125 40675 9183 40681
rect 6779 40477 6837 40483
rect 6779 40474 6791 40477
rect 6748 40452 6791 40474
rect 6730 40400 6736 40452
rect 6788 40443 6791 40452
rect 6825 40443 6837 40477
rect 7742 40468 7748 40520
rect 7800 40508 7806 40520
rect 7929 40511 7987 40517
rect 7929 40508 7941 40511
rect 7800 40480 7941 40508
rect 7800 40468 7806 40480
rect 7929 40477 7941 40480
rect 7975 40477 7987 40511
rect 7929 40471 7987 40477
rect 9217 40511 9275 40517
rect 9217 40477 9229 40511
rect 9263 40508 9275 40511
rect 9674 40508 9680 40520
rect 9263 40480 9680 40508
rect 9263 40477 9275 40480
rect 9217 40471 9275 40477
rect 9674 40468 9680 40480
rect 9732 40468 9738 40520
rect 12618 40468 12624 40520
rect 12676 40508 12682 40520
rect 12713 40511 12771 40517
rect 12713 40508 12725 40511
rect 12676 40480 12725 40508
rect 12676 40468 12682 40480
rect 12713 40477 12725 40480
rect 12759 40477 12771 40511
rect 12713 40471 12771 40477
rect 14734 40468 14740 40520
rect 14792 40508 14798 40520
rect 15565 40511 15623 40517
rect 15565 40508 15577 40511
rect 14792 40480 15577 40508
rect 14792 40468 14798 40480
rect 15565 40477 15577 40480
rect 15611 40508 15623 40511
rect 16025 40511 16083 40517
rect 16025 40508 16037 40511
rect 15611 40480 16037 40508
rect 15611 40477 15623 40480
rect 15565 40471 15623 40477
rect 16025 40477 16037 40480
rect 16071 40477 16083 40511
rect 16025 40471 16083 40477
rect 16114 40468 16120 40520
rect 16172 40508 16178 40520
rect 16281 40511 16339 40517
rect 16281 40508 16293 40511
rect 16172 40480 16293 40508
rect 16172 40468 16178 40480
rect 16281 40477 16293 40480
rect 16327 40477 16339 40511
rect 16281 40471 16339 40477
rect 6788 40437 6837 40443
rect 7009 40443 7067 40449
rect 6788 40400 6794 40437
rect 7009 40409 7021 40443
rect 7055 40409 7067 40443
rect 7009 40403 7067 40409
rect 8113 40443 8171 40449
rect 8113 40409 8125 40443
rect 8159 40440 8171 40443
rect 8294 40440 8300 40452
rect 8159 40412 8300 40440
rect 8159 40409 8171 40412
rect 8113 40403 8171 40409
rect 6454 40332 6460 40384
rect 6512 40372 6518 40384
rect 6641 40375 6699 40381
rect 6641 40372 6653 40375
rect 6512 40344 6653 40372
rect 6512 40332 6518 40344
rect 6641 40341 6653 40344
rect 6687 40341 6699 40375
rect 7024 40372 7052 40403
rect 8294 40400 8300 40412
rect 8352 40400 8358 40452
rect 15320 40443 15378 40449
rect 15320 40409 15332 40443
rect 15366 40440 15378 40443
rect 15470 40440 15476 40452
rect 15366 40412 15476 40440
rect 15366 40409 15378 40412
rect 15320 40403 15378 40409
rect 15470 40400 15476 40412
rect 15528 40400 15534 40452
rect 7926 40372 7932 40384
rect 7024 40344 7932 40372
rect 6641 40335 6699 40341
rect 7926 40332 7932 40344
rect 7984 40332 7990 40384
rect 12710 40332 12716 40384
rect 12768 40372 12774 40384
rect 12897 40375 12955 40381
rect 12897 40372 12909 40375
rect 12768 40344 12909 40372
rect 12768 40332 12774 40344
rect 12897 40341 12909 40344
rect 12943 40341 12955 40375
rect 12897 40335 12955 40341
rect 14185 40375 14243 40381
rect 14185 40341 14197 40375
rect 14231 40372 14243 40375
rect 14642 40372 14648 40384
rect 14231 40344 14648 40372
rect 14231 40341 14243 40344
rect 14185 40335 14243 40341
rect 14642 40332 14648 40344
rect 14700 40332 14706 40384
rect 17402 40372 17408 40384
rect 17363 40344 17408 40372
rect 17402 40332 17408 40344
rect 17460 40332 17466 40384
rect 1104 40282 18860 40304
rect 1104 40230 6880 40282
rect 6932 40230 6944 40282
rect 6996 40230 7008 40282
rect 7060 40230 7072 40282
rect 7124 40230 7136 40282
rect 7188 40230 12811 40282
rect 12863 40230 12875 40282
rect 12927 40230 12939 40282
rect 12991 40230 13003 40282
rect 13055 40230 13067 40282
rect 13119 40230 18860 40282
rect 1104 40208 18860 40230
rect 7561 40171 7619 40177
rect 7561 40137 7573 40171
rect 7607 40168 7619 40171
rect 8110 40168 8116 40180
rect 7607 40140 8116 40168
rect 7607 40137 7619 40140
rect 7561 40131 7619 40137
rect 8110 40128 8116 40140
rect 8168 40128 8174 40180
rect 7837 40103 7895 40109
rect 7837 40069 7849 40103
rect 7883 40100 7895 40103
rect 8018 40100 8024 40112
rect 7883 40072 8024 40100
rect 7883 40069 7895 40072
rect 7837 40063 7895 40069
rect 8018 40060 8024 40072
rect 8076 40060 8082 40112
rect 8754 40100 8760 40112
rect 8128 40072 8760 40100
rect 5626 40032 5632 40044
rect 5587 40004 5632 40032
rect 5626 39992 5632 40004
rect 5684 39992 5690 40044
rect 5825 40035 5883 40041
rect 5825 40001 5837 40035
rect 5871 40032 5883 40035
rect 6546 40032 6552 40044
rect 5871 40004 5948 40032
rect 6507 40004 6552 40032
rect 5871 40001 5883 40004
rect 5825 39995 5883 40001
rect 5920 39964 5948 40004
rect 6546 39992 6552 40004
rect 6604 39992 6610 40044
rect 6638 39992 6644 40044
rect 6696 40032 6702 40044
rect 7742 40041 7748 40044
rect 7720 40035 7748 40041
rect 6696 40004 6868 40032
rect 6696 39992 6702 40004
rect 6840 39976 6868 40004
rect 7720 40001 7732 40035
rect 7720 39995 7748 40001
rect 7742 39992 7748 39995
rect 7800 39992 7806 40044
rect 7926 40032 7932 40044
rect 7887 40004 7932 40032
rect 7926 39992 7932 40004
rect 7984 39992 7990 40044
rect 8128 40041 8156 40072
rect 8754 40060 8760 40072
rect 8812 40060 8818 40112
rect 12710 40060 12716 40112
rect 12768 40100 12774 40112
rect 12866 40103 12924 40109
rect 12866 40100 12878 40103
rect 12768 40072 12878 40100
rect 12768 40060 12774 40072
rect 12866 40069 12878 40072
rect 12912 40069 12924 40103
rect 12866 40063 12924 40069
rect 15378 40060 15384 40112
rect 15436 40100 15442 40112
rect 15436 40072 16574 40100
rect 15436 40060 15442 40072
rect 8112 40035 8170 40041
rect 8112 40001 8124 40035
rect 8158 40001 8170 40035
rect 8112 39995 8170 40001
rect 8205 40035 8263 40041
rect 8205 40001 8217 40035
rect 8251 40032 8263 40035
rect 8938 40032 8944 40044
rect 8251 40004 8944 40032
rect 8251 40001 8263 40004
rect 8205 39995 8263 40001
rect 8938 39992 8944 40004
rect 8996 39992 9002 40044
rect 10226 39992 10232 40044
rect 10284 40032 10290 40044
rect 10505 40035 10563 40041
rect 10505 40032 10517 40035
rect 10284 40004 10517 40032
rect 10284 39992 10290 40004
rect 10505 40001 10517 40004
rect 10551 40001 10563 40035
rect 10505 39995 10563 40001
rect 11977 40035 12035 40041
rect 11977 40001 11989 40035
rect 12023 40032 12035 40035
rect 12066 40032 12072 40044
rect 12023 40004 12072 40032
rect 12023 40001 12035 40004
rect 11977 39995 12035 40001
rect 12066 39992 12072 40004
rect 12124 39992 12130 40044
rect 12161 40035 12219 40041
rect 12161 40001 12173 40035
rect 12207 40032 12219 40035
rect 12526 40032 12532 40044
rect 12207 40004 12532 40032
rect 12207 40001 12219 40004
rect 12161 39995 12219 40001
rect 12526 39992 12532 40004
rect 12584 39992 12590 40044
rect 15004 40035 15062 40041
rect 15004 40001 15016 40035
rect 15050 40032 15062 40035
rect 15562 40032 15568 40044
rect 15050 40004 15568 40032
rect 15050 40001 15062 40004
rect 15004 39995 15062 40001
rect 15562 39992 15568 40004
rect 15620 39992 15626 40044
rect 16546 40032 16574 40072
rect 16853 40035 16911 40041
rect 16853 40032 16865 40035
rect 16546 40004 16865 40032
rect 16853 40001 16865 40004
rect 16899 40001 16911 40035
rect 16853 39995 16911 40001
rect 5994 39964 6000 39976
rect 5907 39936 6000 39964
rect 5994 39924 6000 39936
rect 6052 39964 6058 39976
rect 6730 39964 6736 39976
rect 6052 39936 6736 39964
rect 6052 39924 6058 39936
rect 6730 39924 6736 39936
rect 6788 39924 6794 39976
rect 6822 39924 6828 39976
rect 6880 39964 6886 39976
rect 6880 39936 6925 39964
rect 6880 39924 6886 39936
rect 10318 39924 10324 39976
rect 10376 39964 10382 39976
rect 10413 39967 10471 39973
rect 10413 39964 10425 39967
rect 10376 39936 10425 39964
rect 10376 39924 10382 39936
rect 10413 39933 10425 39936
rect 10459 39933 10471 39967
rect 10413 39927 10471 39933
rect 12621 39967 12679 39973
rect 12621 39933 12633 39967
rect 12667 39933 12679 39967
rect 12621 39927 12679 39933
rect 5534 39788 5540 39840
rect 5592 39828 5598 39840
rect 5813 39831 5871 39837
rect 5813 39828 5825 39831
rect 5592 39800 5825 39828
rect 5592 39788 5598 39800
rect 5813 39797 5825 39800
rect 5859 39797 5871 39831
rect 5813 39791 5871 39797
rect 5902 39788 5908 39840
rect 5960 39828 5966 39840
rect 6748 39837 6776 39924
rect 6365 39831 6423 39837
rect 6365 39828 6377 39831
rect 5960 39800 6377 39828
rect 5960 39788 5966 39800
rect 6365 39797 6377 39800
rect 6411 39797 6423 39831
rect 6365 39791 6423 39797
rect 6733 39831 6791 39837
rect 6733 39797 6745 39831
rect 6779 39828 6791 39831
rect 8110 39828 8116 39840
rect 6779 39800 8116 39828
rect 6779 39797 6791 39800
rect 6733 39791 6791 39797
rect 8110 39788 8116 39800
rect 8168 39788 8174 39840
rect 10778 39828 10784 39840
rect 10739 39800 10784 39828
rect 10778 39788 10784 39800
rect 10836 39788 10842 39840
rect 11698 39788 11704 39840
rect 11756 39828 11762 39840
rect 12069 39831 12127 39837
rect 12069 39828 12081 39831
rect 11756 39800 12081 39828
rect 11756 39788 11762 39800
rect 12069 39797 12081 39800
rect 12115 39797 12127 39831
rect 12636 39828 12664 39927
rect 13814 39924 13820 39976
rect 13872 39964 13878 39976
rect 14734 39964 14740 39976
rect 13872 39936 14740 39964
rect 13872 39924 13878 39936
rect 14734 39924 14740 39936
rect 14792 39924 14798 39976
rect 16666 39924 16672 39976
rect 16724 39964 16730 39976
rect 17037 39967 17095 39973
rect 16724 39936 16769 39964
rect 16724 39924 16730 39936
rect 17037 39933 17049 39967
rect 17083 39933 17095 39967
rect 17037 39927 17095 39933
rect 16114 39896 16120 39908
rect 16027 39868 16120 39896
rect 16114 39856 16120 39868
rect 16172 39896 16178 39908
rect 17052 39896 17080 39927
rect 16172 39868 17080 39896
rect 16172 39856 16178 39868
rect 13814 39828 13820 39840
rect 12636 39800 13820 39828
rect 12069 39791 12127 39797
rect 13814 39788 13820 39800
rect 13872 39788 13878 39840
rect 14001 39831 14059 39837
rect 14001 39797 14013 39831
rect 14047 39828 14059 39831
rect 14458 39828 14464 39840
rect 14047 39800 14464 39828
rect 14047 39797 14059 39800
rect 14001 39791 14059 39797
rect 14458 39788 14464 39800
rect 14516 39828 14522 39840
rect 15102 39828 15108 39840
rect 14516 39800 15108 39828
rect 14516 39788 14522 39800
rect 15102 39788 15108 39800
rect 15160 39788 15166 39840
rect 1104 39738 18860 39760
rect 1104 39686 3915 39738
rect 3967 39686 3979 39738
rect 4031 39686 4043 39738
rect 4095 39686 4107 39738
rect 4159 39686 4171 39738
rect 4223 39686 9846 39738
rect 9898 39686 9910 39738
rect 9962 39686 9974 39738
rect 10026 39686 10038 39738
rect 10090 39686 10102 39738
rect 10154 39686 15776 39738
rect 15828 39686 15840 39738
rect 15892 39686 15904 39738
rect 15956 39686 15968 39738
rect 16020 39686 16032 39738
rect 16084 39686 18860 39738
rect 1104 39664 18860 39686
rect 9674 39584 9680 39636
rect 9732 39624 9738 39636
rect 10781 39627 10839 39633
rect 10781 39624 10793 39627
rect 9732 39596 10793 39624
rect 9732 39584 9738 39596
rect 10781 39593 10793 39596
rect 10827 39593 10839 39627
rect 11882 39624 11888 39636
rect 11843 39596 11888 39624
rect 10781 39587 10839 39593
rect 11882 39584 11888 39596
rect 11940 39584 11946 39636
rect 12618 39584 12624 39636
rect 12676 39624 12682 39636
rect 12805 39627 12863 39633
rect 12805 39624 12817 39627
rect 12676 39596 12817 39624
rect 12676 39584 12682 39596
rect 12805 39593 12817 39596
rect 12851 39593 12863 39627
rect 12805 39587 12863 39593
rect 14737 39627 14795 39633
rect 14737 39593 14749 39627
rect 14783 39624 14795 39627
rect 15102 39624 15108 39636
rect 14783 39596 15108 39624
rect 14783 39593 14795 39596
rect 14737 39587 14795 39593
rect 15102 39584 15108 39596
rect 15160 39584 15166 39636
rect 15378 39584 15384 39636
rect 15436 39624 15442 39636
rect 15436 39596 15608 39624
rect 15436 39584 15442 39596
rect 6365 39559 6423 39565
rect 6365 39525 6377 39559
rect 6411 39525 6423 39559
rect 6365 39519 6423 39525
rect 6380 39488 6408 39519
rect 7558 39516 7564 39568
rect 7616 39556 7622 39568
rect 8389 39559 8447 39565
rect 8389 39556 8401 39559
rect 7616 39528 8401 39556
rect 7616 39516 7622 39528
rect 8389 39525 8401 39528
rect 8435 39525 8447 39559
rect 10226 39556 10232 39568
rect 10187 39528 10232 39556
rect 8389 39519 8447 39525
rect 10226 39516 10232 39528
rect 10284 39516 10290 39568
rect 11054 39556 11060 39568
rect 10967 39528 11060 39556
rect 6825 39491 6883 39497
rect 6825 39488 6837 39491
rect 6380 39460 6837 39488
rect 6825 39457 6837 39460
rect 6871 39488 6883 39491
rect 7374 39488 7380 39500
rect 6871 39460 7380 39488
rect 6871 39457 6883 39460
rect 6825 39451 6883 39457
rect 7374 39448 7380 39460
rect 7432 39448 7438 39500
rect 9950 39488 9956 39500
rect 9911 39460 9956 39488
rect 9950 39448 9956 39460
rect 10008 39448 10014 39500
rect 10980 39497 11008 39528
rect 11054 39516 11060 39528
rect 11112 39556 11118 39568
rect 12250 39556 12256 39568
rect 11112 39528 12256 39556
rect 11112 39516 11118 39528
rect 12250 39516 12256 39528
rect 12308 39516 12314 39568
rect 12636 39528 15516 39556
rect 10965 39491 11023 39497
rect 10965 39457 10977 39491
rect 11011 39457 11023 39491
rect 10965 39451 11023 39457
rect 11977 39491 12035 39497
rect 11977 39457 11989 39491
rect 12023 39488 12035 39491
rect 12526 39488 12532 39500
rect 12023 39460 12532 39488
rect 12023 39457 12035 39460
rect 11977 39451 12035 39457
rect 12526 39448 12532 39460
rect 12584 39448 12590 39500
rect 3602 39380 3608 39432
rect 3660 39420 3666 39432
rect 4985 39423 5043 39429
rect 4985 39420 4997 39423
rect 3660 39392 4997 39420
rect 3660 39380 3666 39392
rect 4985 39389 4997 39392
rect 5031 39420 5043 39423
rect 6362 39420 6368 39432
rect 5031 39392 6368 39420
rect 5031 39389 5043 39392
rect 4985 39383 5043 39389
rect 6362 39380 6368 39392
rect 6420 39380 6426 39432
rect 7101 39423 7159 39429
rect 7101 39389 7113 39423
rect 7147 39389 7159 39423
rect 8110 39420 8116 39432
rect 8071 39392 8116 39420
rect 7101 39383 7159 39389
rect 5252 39355 5310 39361
rect 5252 39321 5264 39355
rect 5298 39352 5310 39355
rect 5902 39352 5908 39364
rect 5298 39324 5908 39352
rect 5298 39321 5310 39324
rect 5252 39315 5310 39321
rect 5902 39312 5908 39324
rect 5960 39312 5966 39364
rect 6822 39312 6828 39364
rect 6880 39312 6886 39364
rect 5718 39244 5724 39296
rect 5776 39284 5782 39296
rect 6840 39284 6868 39312
rect 7116 39284 7144 39383
rect 8110 39380 8116 39392
rect 8168 39380 8174 39432
rect 9861 39423 9919 39429
rect 9861 39389 9873 39423
rect 9907 39420 9919 39423
rect 10689 39423 10747 39429
rect 10689 39420 10701 39423
rect 9907 39392 10701 39420
rect 9907 39389 9919 39392
rect 9861 39383 9919 39389
rect 10689 39389 10701 39392
rect 10735 39389 10747 39423
rect 11698 39420 11704 39432
rect 11659 39392 11704 39420
rect 10689 39383 10747 39389
rect 7926 39312 7932 39364
rect 7984 39352 7990 39364
rect 8389 39355 8447 39361
rect 8389 39352 8401 39355
rect 7984 39324 8401 39352
rect 7984 39312 7990 39324
rect 8389 39321 8401 39324
rect 8435 39321 8447 39355
rect 8389 39315 8447 39321
rect 9766 39312 9772 39364
rect 9824 39352 9830 39364
rect 9876 39352 9904 39383
rect 11698 39380 11704 39392
rect 11756 39380 11762 39432
rect 11790 39380 11796 39432
rect 11848 39420 11854 39432
rect 12636 39429 12664 39528
rect 14553 39491 14611 39497
rect 14553 39457 14565 39491
rect 14599 39488 14611 39491
rect 15194 39488 15200 39500
rect 14599 39460 15200 39488
rect 14599 39457 14611 39460
rect 14553 39451 14611 39457
rect 15194 39448 15200 39460
rect 15252 39448 15258 39500
rect 12437 39423 12495 39429
rect 11848 39392 11893 39420
rect 11848 39380 11854 39392
rect 12437 39389 12449 39423
rect 12483 39389 12495 39423
rect 12437 39383 12495 39389
rect 12621 39423 12679 39429
rect 12621 39389 12633 39423
rect 12667 39389 12679 39423
rect 12621 39383 12679 39389
rect 13541 39423 13599 39429
rect 13541 39389 13553 39423
rect 13587 39420 13599 39423
rect 13587 39392 14596 39420
rect 13587 39389 13599 39392
rect 13541 39383 13599 39389
rect 9824 39324 9904 39352
rect 12452 39352 12480 39383
rect 13446 39352 13452 39364
rect 12452 39324 13452 39352
rect 9824 39312 9830 39324
rect 13446 39312 13452 39324
rect 13504 39312 13510 39364
rect 14182 39312 14188 39364
rect 14240 39352 14246 39364
rect 14461 39355 14519 39361
rect 14461 39352 14473 39355
rect 14240 39324 14473 39352
rect 14240 39312 14246 39324
rect 14461 39321 14473 39324
rect 14507 39321 14519 39355
rect 14568 39352 14596 39392
rect 14642 39380 14648 39432
rect 14700 39420 14706 39432
rect 14737 39423 14795 39429
rect 14737 39420 14749 39423
rect 14700 39392 14749 39420
rect 14700 39380 14706 39392
rect 14737 39389 14749 39392
rect 14783 39389 14795 39423
rect 14737 39383 14795 39389
rect 15381 39355 15439 39361
rect 15381 39352 15393 39355
rect 14568 39324 15393 39352
rect 14461 39315 14519 39321
rect 15381 39321 15393 39324
rect 15427 39321 15439 39355
rect 15488 39352 15516 39528
rect 15580 39488 15608 39596
rect 15746 39516 15752 39568
rect 15804 39556 15810 39568
rect 15804 39528 16528 39556
rect 15804 39516 15810 39528
rect 15580 39460 16436 39488
rect 15580 39429 15608 39460
rect 15565 39423 15623 39429
rect 15565 39389 15577 39423
rect 15611 39389 15623 39423
rect 15565 39383 15623 39389
rect 15654 39380 15660 39432
rect 15712 39420 15718 39432
rect 16408 39429 16436 39460
rect 16500 39429 16528 39528
rect 16393 39423 16451 39429
rect 15712 39392 15757 39420
rect 15712 39380 15718 39392
rect 16393 39389 16405 39423
rect 16439 39389 16451 39423
rect 16393 39383 16451 39389
rect 16485 39423 16543 39429
rect 16485 39389 16497 39423
rect 16531 39389 16543 39423
rect 16485 39383 16543 39389
rect 17954 39352 17960 39364
rect 15488 39324 17960 39352
rect 15381 39315 15439 39321
rect 17954 39312 17960 39324
rect 18012 39312 18018 39364
rect 8205 39287 8263 39293
rect 8205 39284 8217 39287
rect 5776 39256 8217 39284
rect 5776 39244 5782 39256
rect 8205 39253 8217 39256
rect 8251 39284 8263 39287
rect 8478 39284 8484 39296
rect 8251 39256 8484 39284
rect 8251 39253 8263 39256
rect 8205 39247 8263 39253
rect 8478 39244 8484 39256
rect 8536 39244 8542 39296
rect 10410 39244 10416 39296
rect 10468 39284 10474 39296
rect 10965 39287 11023 39293
rect 10965 39284 10977 39287
rect 10468 39256 10977 39284
rect 10468 39244 10474 39256
rect 10965 39253 10977 39256
rect 11011 39253 11023 39287
rect 10965 39247 11023 39253
rect 13170 39244 13176 39296
rect 13228 39284 13234 39296
rect 13357 39287 13415 39293
rect 13357 39284 13369 39287
rect 13228 39256 13369 39284
rect 13228 39244 13234 39256
rect 13357 39253 13369 39256
rect 13403 39253 13415 39287
rect 14918 39284 14924 39296
rect 14879 39256 14924 39284
rect 13357 39247 13415 39253
rect 14918 39244 14924 39256
rect 14976 39244 14982 39296
rect 15930 39244 15936 39296
rect 15988 39284 15994 39296
rect 16209 39287 16267 39293
rect 16209 39284 16221 39287
rect 15988 39256 16221 39284
rect 15988 39244 15994 39256
rect 16209 39253 16221 39256
rect 16255 39253 16267 39287
rect 16209 39247 16267 39253
rect 1104 39194 18860 39216
rect 1104 39142 6880 39194
rect 6932 39142 6944 39194
rect 6996 39142 7008 39194
rect 7060 39142 7072 39194
rect 7124 39142 7136 39194
rect 7188 39142 12811 39194
rect 12863 39142 12875 39194
rect 12927 39142 12939 39194
rect 12991 39142 13003 39194
rect 13055 39142 13067 39194
rect 13119 39142 18860 39194
rect 1104 39120 18860 39142
rect 5635 39083 5693 39089
rect 5635 39049 5647 39083
rect 5681 39080 5693 39083
rect 6546 39080 6552 39092
rect 5681 39052 6552 39080
rect 5681 39049 5693 39052
rect 5635 39043 5693 39049
rect 6546 39040 6552 39052
rect 6604 39040 6610 39092
rect 7745 39083 7803 39089
rect 7745 39049 7757 39083
rect 7791 39080 7803 39083
rect 7926 39080 7932 39092
rect 7791 39052 7932 39080
rect 7791 39049 7803 39052
rect 7745 39043 7803 39049
rect 7926 39040 7932 39052
rect 7984 39040 7990 39092
rect 8938 39080 8944 39092
rect 8899 39052 8944 39080
rect 8938 39040 8944 39052
rect 8996 39040 9002 39092
rect 11054 39080 11060 39092
rect 9692 39052 11060 39080
rect 6362 38972 6368 39024
rect 6420 39012 6426 39024
rect 7282 39012 7288 39024
rect 6420 38984 7288 39012
rect 6420 38972 6426 38984
rect 7282 38972 7288 38984
rect 7340 38972 7346 39024
rect 7944 39012 7972 39040
rect 9692 39012 9720 39052
rect 11054 39040 11060 39052
rect 11112 39040 11118 39092
rect 12066 39080 12072 39092
rect 12027 39052 12072 39080
rect 12066 39040 12072 39052
rect 12124 39040 12130 39092
rect 15102 39080 15108 39092
rect 15063 39052 15108 39080
rect 15102 39040 15108 39052
rect 15160 39040 15166 39092
rect 15562 39040 15568 39092
rect 15620 39080 15626 39092
rect 15749 39083 15807 39089
rect 15749 39080 15761 39083
rect 15620 39052 15761 39080
rect 15620 39040 15626 39052
rect 15749 39049 15761 39052
rect 15795 39049 15807 39083
rect 15749 39043 15807 39049
rect 7944 38984 8616 39012
rect 3602 38944 3608 38956
rect 3563 38916 3608 38944
rect 3602 38904 3608 38916
rect 3660 38904 3666 38956
rect 3694 38904 3700 38956
rect 3752 38944 3758 38956
rect 3861 38947 3919 38953
rect 3861 38944 3873 38947
rect 3752 38916 3873 38944
rect 3752 38904 3758 38916
rect 3861 38913 3873 38916
rect 3907 38913 3919 38947
rect 3861 38907 3919 38913
rect 5537 38947 5595 38953
rect 5537 38913 5549 38947
rect 5583 38913 5595 38947
rect 5718 38944 5724 38956
rect 5679 38916 5724 38944
rect 5537 38907 5595 38913
rect 5552 38876 5580 38907
rect 5718 38904 5724 38916
rect 5776 38904 5782 38956
rect 5813 38947 5871 38953
rect 5813 38913 5825 38947
rect 5859 38944 5871 38947
rect 5994 38944 6000 38956
rect 5859 38916 6000 38944
rect 5859 38913 5871 38916
rect 5813 38907 5871 38913
rect 5994 38904 6000 38916
rect 6052 38904 6058 38956
rect 6638 38953 6644 38956
rect 6632 38907 6644 38953
rect 6696 38944 6702 38956
rect 8202 38944 8208 38956
rect 6696 38916 6732 38944
rect 8163 38916 8208 38944
rect 6638 38904 6644 38907
rect 6696 38904 6702 38916
rect 8202 38904 8208 38916
rect 8260 38904 8266 38956
rect 8386 38944 8392 38956
rect 8347 38916 8392 38944
rect 8386 38904 8392 38916
rect 8444 38904 8450 38956
rect 8588 38953 8616 38984
rect 9600 38984 9720 39012
rect 9861 39015 9919 39021
rect 8573 38947 8631 38953
rect 8573 38913 8585 38947
rect 8619 38913 8631 38947
rect 8754 38944 8760 38956
rect 8715 38916 8760 38944
rect 8573 38907 8631 38913
rect 8754 38904 8760 38916
rect 8812 38904 8818 38956
rect 9600 38953 9628 38984
rect 9861 38981 9873 39015
rect 9907 39012 9919 39015
rect 10502 39012 10508 39024
rect 9907 38984 10508 39012
rect 9907 38981 9919 38984
rect 9861 38975 9919 38981
rect 10502 38972 10508 38984
rect 10560 38972 10566 39024
rect 11885 39015 11943 39021
rect 11885 38981 11897 39015
rect 11931 39012 11943 39015
rect 12434 39012 12440 39024
rect 11931 38984 12440 39012
rect 11931 38981 11943 38984
rect 11885 38975 11943 38981
rect 12434 38972 12440 38984
rect 12492 38972 12498 39024
rect 13814 39012 13820 39024
rect 12912 38984 13820 39012
rect 9585 38947 9643 38953
rect 9585 38913 9597 38947
rect 9631 38913 9643 38947
rect 9585 38907 9643 38913
rect 9674 38904 9680 38956
rect 9732 38944 9738 38956
rect 10410 38944 10416 38956
rect 9732 38916 9777 38944
rect 10371 38916 10416 38944
rect 9732 38904 9738 38916
rect 10410 38904 10416 38916
rect 10468 38904 10474 38956
rect 10689 38947 10747 38953
rect 10689 38913 10701 38947
rect 10735 38944 10747 38947
rect 11701 38947 11759 38953
rect 10735 38916 10824 38944
rect 10735 38913 10747 38916
rect 10689 38907 10747 38913
rect 6362 38876 6368 38888
rect 5552 38848 5672 38876
rect 6323 38848 6368 38876
rect 4522 38700 4528 38752
rect 4580 38740 4586 38752
rect 4985 38743 5043 38749
rect 4985 38740 4997 38743
rect 4580 38712 4997 38740
rect 4580 38700 4586 38712
rect 4985 38709 4997 38712
rect 5031 38709 5043 38743
rect 5644 38740 5672 38848
rect 6362 38836 6368 38848
rect 6420 38836 6426 38888
rect 8018 38836 8024 38888
rect 8076 38876 8082 38888
rect 8481 38879 8539 38885
rect 8481 38876 8493 38879
rect 8076 38848 8493 38876
rect 8076 38836 8082 38848
rect 8481 38845 8493 38848
rect 8527 38845 8539 38879
rect 8481 38839 8539 38845
rect 10226 38836 10232 38888
rect 10284 38876 10290 38888
rect 10505 38879 10563 38885
rect 10505 38876 10517 38879
rect 10284 38848 10517 38876
rect 10284 38836 10290 38848
rect 10505 38845 10517 38848
rect 10551 38845 10563 38879
rect 10505 38839 10563 38845
rect 9861 38811 9919 38817
rect 9861 38777 9873 38811
rect 9907 38808 9919 38811
rect 10318 38808 10324 38820
rect 9907 38780 10324 38808
rect 9907 38777 9919 38780
rect 9861 38771 9919 38777
rect 10318 38768 10324 38780
rect 10376 38768 10382 38820
rect 10594 38808 10600 38820
rect 10555 38780 10600 38808
rect 10594 38768 10600 38780
rect 10652 38768 10658 38820
rect 10796 38808 10824 38916
rect 11701 38913 11713 38947
rect 11747 38944 11759 38947
rect 12250 38944 12256 38956
rect 11747 38916 12256 38944
rect 11747 38913 11759 38916
rect 11701 38907 11759 38913
rect 12250 38904 12256 38916
rect 12308 38904 12314 38956
rect 12912 38953 12940 38984
rect 13814 38972 13820 38984
rect 13872 38972 13878 39024
rect 14642 38972 14648 39024
rect 14700 39012 14706 39024
rect 15289 39015 15347 39021
rect 15289 39012 15301 39015
rect 14700 38984 15301 39012
rect 14700 38972 14706 38984
rect 15289 38981 15301 38984
rect 15335 39012 15347 39015
rect 15654 39012 15660 39024
rect 15335 38984 15660 39012
rect 15335 38981 15347 38984
rect 15289 38975 15347 38981
rect 15654 38972 15660 38984
rect 15712 38972 15718 39024
rect 13170 38953 13176 38956
rect 12897 38947 12955 38953
rect 12897 38913 12909 38947
rect 12943 38913 12955 38947
rect 13164 38944 13176 38953
rect 13131 38916 13176 38944
rect 12897 38907 12955 38913
rect 13164 38907 13176 38916
rect 13170 38904 13176 38907
rect 13228 38904 13234 38956
rect 14182 38904 14188 38956
rect 14240 38944 14246 38956
rect 14921 38947 14979 38953
rect 14921 38944 14933 38947
rect 14240 38916 14933 38944
rect 14240 38904 14246 38916
rect 14921 38913 14933 38916
rect 14967 38913 14979 38947
rect 14921 38907 14979 38913
rect 15013 38947 15071 38953
rect 15013 38913 15025 38947
rect 15059 38944 15071 38947
rect 15194 38944 15200 38956
rect 15059 38916 15200 38944
rect 15059 38913 15071 38916
rect 15013 38907 15071 38913
rect 15194 38904 15200 38916
rect 15252 38944 15258 38956
rect 15746 38944 15752 38956
rect 15252 38916 15752 38944
rect 15252 38904 15258 38916
rect 15746 38904 15752 38916
rect 15804 38904 15810 38956
rect 15930 38944 15936 38956
rect 15891 38916 15936 38944
rect 15930 38904 15936 38916
rect 15988 38904 15994 38956
rect 10873 38879 10931 38885
rect 10873 38845 10885 38879
rect 10919 38876 10931 38879
rect 11790 38876 11796 38888
rect 10919 38848 11796 38876
rect 10919 38845 10931 38848
rect 10873 38839 10931 38845
rect 11790 38836 11796 38848
rect 11848 38836 11854 38888
rect 10962 38808 10968 38820
rect 10796 38780 10968 38808
rect 10962 38768 10968 38780
rect 11020 38768 11026 38820
rect 7834 38740 7840 38752
rect 5644 38712 7840 38740
rect 4985 38703 5043 38709
rect 7834 38700 7840 38712
rect 7892 38700 7898 38752
rect 14182 38700 14188 38752
rect 14240 38740 14246 38752
rect 14277 38743 14335 38749
rect 14277 38740 14289 38743
rect 14240 38712 14289 38740
rect 14240 38700 14246 38712
rect 14277 38709 14289 38712
rect 14323 38709 14335 38743
rect 14277 38703 14335 38709
rect 14366 38700 14372 38752
rect 14424 38740 14430 38752
rect 14737 38743 14795 38749
rect 14737 38740 14749 38743
rect 14424 38712 14749 38740
rect 14424 38700 14430 38712
rect 14737 38709 14749 38712
rect 14783 38709 14795 38743
rect 14737 38703 14795 38709
rect 1104 38650 18860 38672
rect 1104 38598 3915 38650
rect 3967 38598 3979 38650
rect 4031 38598 4043 38650
rect 4095 38598 4107 38650
rect 4159 38598 4171 38650
rect 4223 38598 9846 38650
rect 9898 38598 9910 38650
rect 9962 38598 9974 38650
rect 10026 38598 10038 38650
rect 10090 38598 10102 38650
rect 10154 38598 15776 38650
rect 15828 38598 15840 38650
rect 15892 38598 15904 38650
rect 15956 38598 15968 38650
rect 16020 38598 16032 38650
rect 16084 38598 18860 38650
rect 1104 38576 18860 38598
rect 12526 38536 12532 38548
rect 12487 38508 12532 38536
rect 12526 38496 12532 38508
rect 12584 38496 12590 38548
rect 15194 38496 15200 38548
rect 15252 38536 15258 38548
rect 15473 38539 15531 38545
rect 15473 38536 15485 38539
rect 15252 38508 15485 38536
rect 15252 38496 15258 38508
rect 15473 38505 15485 38508
rect 15519 38505 15531 38539
rect 15473 38499 15531 38505
rect 6641 38471 6699 38477
rect 6641 38437 6653 38471
rect 6687 38468 6699 38471
rect 6730 38468 6736 38480
rect 6687 38440 6736 38468
rect 6687 38437 6699 38440
rect 6641 38431 6699 38437
rect 6730 38428 6736 38440
rect 6788 38468 6794 38480
rect 10965 38471 11023 38477
rect 6788 38440 7144 38468
rect 6788 38428 6794 38440
rect 7116 38409 7144 38440
rect 10965 38437 10977 38471
rect 11011 38468 11023 38471
rect 11054 38468 11060 38480
rect 11011 38440 11060 38468
rect 11011 38437 11023 38440
rect 10965 38431 11023 38437
rect 11054 38428 11060 38440
rect 11112 38428 11118 38480
rect 7101 38403 7159 38409
rect 7101 38369 7113 38403
rect 7147 38369 7159 38403
rect 7101 38363 7159 38369
rect 7377 38403 7435 38409
rect 7377 38369 7389 38403
rect 7423 38400 7435 38403
rect 8110 38400 8116 38412
rect 7423 38372 8116 38400
rect 7423 38369 7435 38372
rect 7377 38363 7435 38369
rect 8110 38360 8116 38372
rect 8168 38360 8174 38412
rect 9766 38400 9772 38412
rect 9727 38372 9772 38400
rect 9766 38360 9772 38372
rect 9824 38400 9830 38412
rect 10318 38400 10324 38412
rect 9824 38372 10324 38400
rect 9824 38360 9830 38372
rect 10318 38360 10324 38372
rect 10376 38400 10382 38412
rect 11701 38403 11759 38409
rect 10376 38372 10824 38400
rect 10376 38360 10382 38372
rect 3786 38332 3792 38344
rect 3747 38304 3792 38332
rect 3786 38292 3792 38304
rect 3844 38292 3850 38344
rect 3973 38335 4031 38341
rect 3973 38301 3985 38335
rect 4019 38332 4031 38335
rect 4890 38332 4896 38344
rect 4019 38304 4896 38332
rect 4019 38301 4031 38304
rect 3973 38295 4031 38301
rect 4890 38292 4896 38304
rect 4948 38292 4954 38344
rect 5261 38335 5319 38341
rect 5261 38301 5273 38335
rect 5307 38332 5319 38335
rect 6362 38332 6368 38344
rect 5307 38304 6368 38332
rect 5307 38301 5319 38304
rect 5261 38295 5319 38301
rect 5644 38276 5672 38304
rect 6362 38292 6368 38304
rect 6420 38292 6426 38344
rect 9674 38292 9680 38344
rect 9732 38332 9738 38344
rect 10226 38332 10232 38344
rect 9732 38304 10232 38332
rect 9732 38292 9738 38304
rect 10226 38292 10232 38304
rect 10284 38292 10290 38344
rect 10796 38341 10824 38372
rect 11701 38369 11713 38403
rect 11747 38400 11759 38403
rect 11790 38400 11796 38412
rect 11747 38372 11796 38400
rect 11747 38369 11759 38372
rect 11701 38363 11759 38369
rect 11790 38360 11796 38372
rect 11848 38360 11854 38412
rect 13814 38360 13820 38412
rect 13872 38400 13878 38412
rect 14093 38403 14151 38409
rect 14093 38400 14105 38403
rect 13872 38372 14105 38400
rect 13872 38360 13878 38372
rect 14093 38369 14105 38372
rect 14139 38369 14151 38403
rect 14093 38363 14151 38369
rect 10781 38335 10839 38341
rect 10781 38301 10793 38335
rect 10827 38301 10839 38335
rect 11606 38332 11612 38344
rect 11567 38304 11612 38332
rect 10781 38295 10839 38301
rect 11606 38292 11612 38304
rect 11664 38292 11670 38344
rect 12250 38292 12256 38344
rect 12308 38332 12314 38344
rect 12437 38335 12495 38341
rect 12437 38332 12449 38335
rect 12308 38304 12449 38332
rect 12308 38292 12314 38304
rect 12437 38301 12449 38304
rect 12483 38301 12495 38335
rect 12437 38295 12495 38301
rect 12526 38292 12532 38344
rect 12584 38332 12590 38344
rect 12621 38335 12679 38341
rect 12621 38332 12633 38335
rect 12584 38304 12633 38332
rect 12584 38292 12590 38304
rect 12621 38301 12633 38304
rect 12667 38301 12679 38335
rect 13354 38332 13360 38344
rect 13315 38304 13360 38332
rect 12621 38295 12679 38301
rect 13354 38292 13360 38304
rect 13412 38292 13418 38344
rect 5534 38273 5540 38276
rect 5528 38264 5540 38273
rect 5495 38236 5540 38264
rect 5528 38227 5540 38236
rect 5534 38224 5540 38227
rect 5592 38224 5598 38276
rect 5626 38224 5632 38276
rect 5684 38224 5690 38276
rect 14338 38267 14396 38273
rect 14338 38264 14350 38267
rect 13556 38236 14350 38264
rect 3973 38199 4031 38205
rect 3973 38165 3985 38199
rect 4019 38196 4031 38199
rect 4246 38196 4252 38208
rect 4019 38168 4252 38196
rect 4019 38165 4031 38168
rect 3973 38159 4031 38165
rect 4246 38156 4252 38168
rect 4304 38156 4310 38208
rect 10045 38199 10103 38205
rect 10045 38165 10057 38199
rect 10091 38196 10103 38199
rect 10594 38196 10600 38208
rect 10091 38168 10600 38196
rect 10091 38165 10103 38168
rect 10045 38159 10103 38165
rect 10594 38156 10600 38168
rect 10652 38156 10658 38208
rect 11977 38199 12035 38205
rect 11977 38165 11989 38199
rect 12023 38196 12035 38199
rect 12250 38196 12256 38208
rect 12023 38168 12256 38196
rect 12023 38165 12035 38168
rect 11977 38159 12035 38165
rect 12250 38156 12256 38168
rect 12308 38156 12314 38208
rect 13556 38205 13584 38236
rect 14338 38233 14350 38236
rect 14384 38233 14396 38267
rect 14338 38227 14396 38233
rect 13541 38199 13599 38205
rect 13541 38165 13553 38199
rect 13587 38165 13599 38199
rect 13541 38159 13599 38165
rect 1104 38106 18860 38128
rect 1104 38054 6880 38106
rect 6932 38054 6944 38106
rect 6996 38054 7008 38106
rect 7060 38054 7072 38106
rect 7124 38054 7136 38106
rect 7188 38054 12811 38106
rect 12863 38054 12875 38106
rect 12927 38054 12939 38106
rect 12991 38054 13003 38106
rect 13055 38054 13067 38106
rect 13119 38054 18860 38106
rect 1104 38032 18860 38054
rect 7377 37995 7435 38001
rect 7377 37961 7389 37995
rect 7423 37992 7435 37995
rect 8202 37992 8208 38004
rect 7423 37964 8208 37992
rect 7423 37961 7435 37964
rect 7377 37955 7435 37961
rect 8202 37952 8208 37964
rect 8260 37952 8266 38004
rect 9674 37952 9680 38004
rect 9732 37952 9738 38004
rect 12526 37952 12532 38004
rect 12584 37992 12590 38004
rect 12897 37995 12955 38001
rect 12897 37992 12909 37995
rect 12584 37964 12909 37992
rect 12584 37952 12590 37964
rect 12897 37961 12909 37964
rect 12943 37961 12955 37995
rect 12897 37955 12955 37961
rect 5626 37924 5632 37936
rect 3896 37896 5632 37924
rect 2774 37816 2780 37868
rect 2832 37856 2838 37868
rect 3896 37865 3924 37896
rect 5626 37884 5632 37896
rect 5684 37884 5690 37936
rect 6730 37884 6736 37936
rect 6788 37924 6794 37936
rect 8113 37927 8171 37933
rect 6788 37896 6960 37924
rect 6788 37884 6794 37896
rect 2869 37859 2927 37865
rect 2869 37856 2881 37859
rect 2832 37828 2881 37856
rect 2832 37816 2838 37828
rect 2869 37825 2881 37828
rect 2915 37825 2927 37859
rect 2869 37819 2927 37825
rect 3881 37859 3939 37865
rect 3881 37825 3893 37859
rect 3927 37825 3939 37859
rect 3881 37819 3939 37825
rect 4148 37859 4206 37865
rect 4148 37825 4160 37859
rect 4194 37856 4206 37859
rect 4706 37856 4712 37868
rect 4194 37828 4712 37856
rect 4194 37825 4206 37828
rect 4148 37819 4206 37825
rect 4706 37816 4712 37828
rect 4764 37816 4770 37868
rect 6546 37816 6552 37868
rect 6604 37856 6610 37868
rect 6932 37865 6960 37896
rect 8113 37893 8125 37927
rect 8159 37924 8171 37927
rect 8754 37924 8760 37936
rect 8159 37896 8760 37924
rect 8159 37893 8171 37896
rect 8113 37887 8171 37893
rect 8754 37884 8760 37896
rect 8812 37884 8818 37936
rect 9705 37871 9733 37952
rect 10686 37884 10692 37936
rect 10744 37924 10750 37936
rect 10870 37924 10876 37936
rect 10744 37896 10876 37924
rect 10744 37884 10750 37896
rect 10870 37884 10876 37896
rect 10928 37884 10934 37936
rect 13814 37924 13820 37936
rect 11532 37896 13820 37924
rect 6825 37859 6883 37865
rect 6825 37856 6837 37859
rect 6604 37828 6837 37856
rect 6604 37816 6610 37828
rect 6825 37825 6837 37828
rect 6871 37825 6883 37859
rect 6825 37819 6883 37825
rect 6917 37859 6975 37865
rect 6917 37825 6929 37859
rect 6963 37825 6975 37859
rect 6917 37819 6975 37825
rect 7101 37859 7159 37865
rect 7101 37825 7113 37859
rect 7147 37825 7159 37859
rect 7101 37819 7159 37825
rect 7193 37859 7251 37865
rect 7193 37825 7205 37859
rect 7239 37856 7251 37859
rect 7374 37856 7380 37868
rect 7239 37828 7380 37856
rect 7239 37825 7251 37828
rect 7193 37819 7251 37825
rect 3142 37788 3148 37800
rect 3103 37760 3148 37788
rect 3142 37748 3148 37760
rect 3200 37748 3206 37800
rect 7116 37788 7144 37819
rect 7374 37816 7380 37828
rect 7432 37816 7438 37868
rect 7742 37816 7748 37868
rect 7800 37856 7806 37868
rect 8205 37859 8263 37865
rect 8205 37856 8217 37859
rect 7800 37828 8217 37856
rect 7800 37816 7806 37828
rect 8205 37825 8217 37828
rect 8251 37825 8263 37859
rect 8846 37856 8852 37868
rect 8807 37828 8852 37856
rect 8205 37819 8263 37825
rect 8846 37816 8852 37828
rect 8904 37816 8910 37868
rect 9674 37865 9733 37871
rect 9585 37859 9643 37865
rect 9585 37825 9597 37859
rect 9631 37825 9643 37859
rect 9674 37831 9686 37865
rect 9720 37834 9733 37865
rect 9720 37831 9732 37834
rect 9674 37825 9732 37831
rect 9585 37819 9643 37825
rect 8018 37788 8024 37800
rect 7116 37760 8024 37788
rect 8018 37748 8024 37760
rect 8076 37748 8082 37800
rect 8294 37748 8300 37800
rect 8352 37788 8358 37800
rect 8757 37791 8815 37797
rect 8757 37788 8769 37791
rect 8352 37760 8769 37788
rect 8352 37748 8358 37760
rect 8757 37757 8769 37760
rect 8803 37757 8815 37791
rect 9600 37788 9628 37819
rect 9766 37816 9772 37868
rect 9824 37865 9830 37868
rect 9824 37856 9832 37865
rect 9953 37859 10011 37865
rect 9824 37828 9869 37856
rect 9824 37819 9832 37828
rect 9953 37825 9965 37859
rect 9999 37856 10011 37859
rect 10594 37856 10600 37868
rect 9999 37828 10364 37856
rect 10555 37828 10600 37856
rect 9999 37825 10011 37828
rect 9953 37819 10011 37825
rect 9824 37816 9830 37819
rect 10226 37788 10232 37800
rect 9600 37760 10232 37788
rect 8757 37751 8815 37757
rect 10226 37748 10232 37760
rect 10284 37748 10290 37800
rect 10336 37788 10364 37828
rect 10594 37816 10600 37828
rect 10652 37816 10658 37868
rect 11532 37865 11560 37896
rect 13814 37884 13820 37896
rect 13872 37884 13878 37936
rect 11790 37865 11796 37868
rect 11517 37859 11575 37865
rect 11517 37825 11529 37859
rect 11563 37825 11575 37859
rect 11517 37819 11575 37825
rect 11784 37819 11796 37865
rect 11848 37856 11854 37868
rect 13998 37856 14004 37868
rect 11848 37828 11884 37856
rect 13959 37828 14004 37856
rect 11790 37816 11796 37819
rect 11848 37816 11854 37828
rect 13998 37816 14004 37828
rect 14056 37816 14062 37868
rect 14182 37856 14188 37868
rect 14143 37828 14188 37856
rect 14182 37816 14188 37828
rect 14240 37816 14246 37868
rect 10686 37788 10692 37800
rect 10336 37760 10692 37788
rect 10686 37748 10692 37760
rect 10744 37748 10750 37800
rect 10781 37791 10839 37797
rect 10781 37757 10793 37791
rect 10827 37788 10839 37791
rect 10962 37788 10968 37800
rect 10827 37760 10968 37788
rect 10827 37757 10839 37760
rect 10781 37751 10839 37757
rect 10962 37748 10968 37760
rect 11020 37748 11026 37800
rect 13354 37748 13360 37800
rect 13412 37788 13418 37800
rect 13817 37791 13875 37797
rect 13817 37788 13829 37791
rect 13412 37760 13829 37788
rect 13412 37748 13418 37760
rect 13817 37757 13829 37760
rect 13863 37757 13875 37791
rect 13817 37751 13875 37757
rect 2958 37652 2964 37664
rect 2919 37624 2964 37652
rect 2958 37612 2964 37624
rect 3016 37612 3022 37664
rect 3053 37655 3111 37661
rect 3053 37621 3065 37655
rect 3099 37652 3111 37655
rect 5074 37652 5080 37664
rect 3099 37624 5080 37652
rect 3099 37621 3111 37624
rect 3053 37615 3111 37621
rect 5074 37612 5080 37624
rect 5132 37612 5138 37664
rect 5261 37655 5319 37661
rect 5261 37621 5273 37655
rect 5307 37652 5319 37655
rect 5350 37652 5356 37664
rect 5307 37624 5356 37652
rect 5307 37621 5319 37624
rect 5261 37615 5319 37621
rect 5350 37612 5356 37624
rect 5408 37612 5414 37664
rect 9309 37655 9367 37661
rect 9309 37621 9321 37655
rect 9355 37652 9367 37655
rect 9398 37652 9404 37664
rect 9355 37624 9404 37652
rect 9355 37621 9367 37624
rect 9309 37615 9367 37621
rect 9398 37612 9404 37624
rect 9456 37612 9462 37664
rect 10410 37652 10416 37664
rect 10371 37624 10416 37652
rect 10410 37612 10416 37624
rect 10468 37612 10474 37664
rect 1104 37562 18860 37584
rect 1104 37510 3915 37562
rect 3967 37510 3979 37562
rect 4031 37510 4043 37562
rect 4095 37510 4107 37562
rect 4159 37510 4171 37562
rect 4223 37510 9846 37562
rect 9898 37510 9910 37562
rect 9962 37510 9974 37562
rect 10026 37510 10038 37562
rect 10090 37510 10102 37562
rect 10154 37510 15776 37562
rect 15828 37510 15840 37562
rect 15892 37510 15904 37562
rect 15956 37510 15968 37562
rect 16020 37510 16032 37562
rect 16084 37510 18860 37562
rect 1104 37488 18860 37510
rect 6638 37448 6644 37460
rect 6599 37420 6644 37448
rect 6638 37408 6644 37420
rect 6696 37408 6702 37460
rect 7193 37451 7251 37457
rect 7193 37417 7205 37451
rect 7239 37448 7251 37451
rect 7282 37448 7288 37460
rect 7239 37420 7288 37448
rect 7239 37417 7251 37420
rect 7193 37411 7251 37417
rect 7282 37408 7288 37420
rect 7340 37408 7346 37460
rect 10410 37448 10416 37460
rect 10371 37420 10416 37448
rect 10410 37408 10416 37420
rect 10468 37408 10474 37460
rect 11790 37448 11796 37460
rect 11751 37420 11796 37448
rect 11790 37408 11796 37420
rect 11848 37408 11854 37460
rect 4890 37380 4896 37392
rect 4172 37352 4896 37380
rect 2225 37247 2283 37253
rect 2225 37213 2237 37247
rect 2271 37213 2283 37247
rect 2225 37207 2283 37213
rect 2409 37247 2467 37253
rect 2409 37213 2421 37247
rect 2455 37244 2467 37247
rect 3142 37244 3148 37256
rect 2455 37216 3148 37244
rect 2455 37213 2467 37216
rect 2409 37207 2467 37213
rect 2240 37176 2268 37207
rect 3142 37204 3148 37216
rect 3200 37204 3206 37256
rect 4172 37253 4200 37352
rect 4890 37340 4896 37352
rect 4948 37340 4954 37392
rect 6549 37383 6607 37389
rect 6549 37349 6561 37383
rect 6595 37380 6607 37383
rect 7558 37380 7564 37392
rect 6595 37352 7564 37380
rect 6595 37349 6607 37352
rect 6549 37343 6607 37349
rect 7558 37340 7564 37352
rect 7616 37340 7622 37392
rect 7926 37340 7932 37392
rect 7984 37380 7990 37392
rect 8202 37380 8208 37392
rect 7984 37352 8208 37380
rect 7984 37340 7990 37352
rect 8202 37340 8208 37352
rect 8260 37340 8266 37392
rect 9766 37340 9772 37392
rect 9824 37380 9830 37392
rect 10321 37383 10379 37389
rect 10321 37380 10333 37383
rect 9824 37352 10333 37380
rect 9824 37340 9830 37352
rect 10321 37349 10333 37352
rect 10367 37349 10379 37383
rect 10870 37380 10876 37392
rect 10321 37343 10379 37349
rect 10428 37352 10876 37380
rect 4982 37312 4988 37324
rect 4943 37284 4988 37312
rect 4982 37272 4988 37284
rect 5040 37272 5046 37324
rect 7466 37272 7472 37324
rect 7524 37312 7530 37324
rect 8941 37315 8999 37321
rect 8941 37312 8953 37315
rect 7524 37284 8953 37312
rect 7524 37272 7530 37284
rect 8941 37281 8953 37284
rect 8987 37281 8999 37315
rect 10229 37315 10287 37321
rect 10229 37312 10241 37315
rect 8941 37275 8999 37281
rect 9140 37284 10241 37312
rect 9140 37256 9168 37284
rect 10229 37281 10241 37284
rect 10275 37312 10287 37315
rect 10428 37312 10456 37352
rect 10870 37340 10876 37352
rect 10928 37340 10934 37392
rect 10275 37284 10456 37312
rect 10275 37281 10287 37284
rect 10229 37275 10287 37281
rect 10686 37272 10692 37324
rect 10744 37312 10750 37324
rect 12345 37315 12403 37321
rect 12345 37312 12357 37315
rect 10744 37284 11100 37312
rect 10744 37272 10750 37284
rect 4065 37247 4123 37253
rect 4065 37213 4077 37247
rect 4111 37213 4123 37247
rect 4065 37207 4123 37213
rect 4157 37247 4215 37253
rect 4157 37213 4169 37247
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 2869 37179 2927 37185
rect 2869 37176 2881 37179
rect 2240 37148 2881 37176
rect 2869 37145 2881 37148
rect 2915 37145 2927 37179
rect 2869 37139 2927 37145
rect 3053 37179 3111 37185
rect 3053 37145 3065 37179
rect 3099 37145 3111 37179
rect 3053 37139 3111 37145
rect 3237 37179 3295 37185
rect 3237 37145 3249 37179
rect 3283 37176 3295 37179
rect 3602 37176 3608 37188
rect 3283 37148 3608 37176
rect 3283 37145 3295 37148
rect 3237 37139 3295 37145
rect 2409 37111 2467 37117
rect 2409 37077 2421 37111
rect 2455 37108 2467 37111
rect 2774 37108 2780 37120
rect 2455 37080 2780 37108
rect 2455 37077 2467 37080
rect 2409 37071 2467 37077
rect 2774 37068 2780 37080
rect 2832 37068 2838 37120
rect 3068 37108 3096 37139
rect 3602 37136 3608 37148
rect 3660 37136 3666 37188
rect 3694 37136 3700 37188
rect 3752 37176 3758 37188
rect 3789 37179 3847 37185
rect 3789 37176 3801 37179
rect 3752 37148 3801 37176
rect 3752 37136 3758 37148
rect 3789 37145 3801 37148
rect 3835 37145 3847 37179
rect 3789 37139 3847 37145
rect 4080 37176 4108 37207
rect 4246 37204 4252 37256
rect 4304 37244 4310 37256
rect 4304 37216 4349 37244
rect 4304 37204 4310 37216
rect 4430 37204 4436 37256
rect 4488 37244 4494 37256
rect 5074 37244 5080 37256
rect 4488 37216 4533 37244
rect 5035 37216 5080 37244
rect 4488 37204 4494 37216
rect 5074 37204 5080 37216
rect 5132 37204 5138 37256
rect 6641 37247 6699 37253
rect 6641 37213 6653 37247
rect 6687 37213 6699 37247
rect 6641 37207 6699 37213
rect 8113 37247 8171 37253
rect 8113 37213 8125 37247
rect 8159 37244 8171 37247
rect 9122 37244 9128 37256
rect 8159 37216 9128 37244
rect 8159 37213 8171 37216
rect 8113 37207 8171 37213
rect 4522 37176 4528 37188
rect 4080 37148 4528 37176
rect 4080 37108 4108 37148
rect 4522 37136 4528 37148
rect 4580 37136 4586 37188
rect 5534 37136 5540 37188
rect 5592 37176 5598 37188
rect 5718 37176 5724 37188
rect 5592 37148 5724 37176
rect 5592 37136 5598 37148
rect 5718 37136 5724 37148
rect 5776 37176 5782 37188
rect 6365 37179 6423 37185
rect 6365 37176 6377 37179
rect 5776 37148 6377 37176
rect 5776 37136 5782 37148
rect 6365 37145 6377 37148
rect 6411 37145 6423 37179
rect 6365 37139 6423 37145
rect 6454 37136 6460 37188
rect 6512 37176 6518 37188
rect 6656 37176 6684 37207
rect 9122 37204 9128 37216
rect 9180 37204 9186 37256
rect 9217 37247 9275 37253
rect 9217 37213 9229 37247
rect 9263 37213 9275 37247
rect 10502 37244 10508 37256
rect 10463 37216 10508 37244
rect 9217 37207 9275 37213
rect 7282 37176 7288 37188
rect 6512 37148 6684 37176
rect 7243 37148 7288 37176
rect 6512 37136 6518 37148
rect 7282 37136 7288 37148
rect 7340 37136 7346 37188
rect 7558 37136 7564 37188
rect 7616 37176 7622 37188
rect 7834 37176 7840 37188
rect 7616 37148 7840 37176
rect 7616 37136 7622 37148
rect 7834 37136 7840 37148
rect 7892 37136 7898 37188
rect 8021 37179 8079 37185
rect 8021 37145 8033 37179
rect 8067 37176 8079 37179
rect 8294 37176 8300 37188
rect 8067 37148 8300 37176
rect 8067 37145 8079 37148
rect 8021 37139 8079 37145
rect 8294 37136 8300 37148
rect 8352 37176 8358 37188
rect 9232 37176 9260 37207
rect 10502 37204 10508 37216
rect 10560 37204 10566 37256
rect 11072 37244 11100 37284
rect 11348 37284 12357 37312
rect 11146 37244 11152 37256
rect 11072 37216 11152 37244
rect 11146 37204 11152 37216
rect 11204 37204 11210 37256
rect 11348 37253 11376 37284
rect 12345 37281 12357 37284
rect 12391 37281 12403 37315
rect 12345 37275 12403 37281
rect 11333 37247 11391 37253
rect 11333 37213 11345 37247
rect 11379 37213 11391 37247
rect 11333 37207 11391 37213
rect 11425 37247 11483 37253
rect 11425 37213 11437 37247
rect 11471 37213 11483 37247
rect 11425 37207 11483 37213
rect 11517 37247 11575 37253
rect 11517 37213 11529 37247
rect 11563 37213 11575 37247
rect 12250 37244 12256 37256
rect 12211 37216 12256 37244
rect 11517 37207 11575 37213
rect 8352 37148 9260 37176
rect 8352 37136 8358 37148
rect 5442 37108 5448 37120
rect 3068 37080 4108 37108
rect 5403 37080 5448 37108
rect 5442 37068 5448 37080
rect 5500 37068 5506 37120
rect 7926 37108 7932 37120
rect 7984 37117 7990 37120
rect 7893 37080 7932 37108
rect 7926 37068 7932 37080
rect 7984 37071 7993 37117
rect 11440 37108 11468 37207
rect 11532 37176 11560 37207
rect 12250 37204 12256 37216
rect 12308 37204 12314 37256
rect 12437 37247 12495 37253
rect 12437 37213 12449 37247
rect 12483 37244 12495 37247
rect 13262 37244 13268 37256
rect 12483 37216 13268 37244
rect 12483 37213 12495 37216
rect 12437 37207 12495 37213
rect 12526 37176 12532 37188
rect 11532 37148 12532 37176
rect 12526 37136 12532 37148
rect 12584 37136 12590 37188
rect 12342 37108 12348 37120
rect 11440 37080 12348 37108
rect 7984 37068 7990 37071
rect 12342 37068 12348 37080
rect 12400 37108 12406 37120
rect 12636 37108 12664 37216
rect 13262 37204 13268 37216
rect 13320 37204 13326 37256
rect 12400 37080 12664 37108
rect 12400 37068 12406 37080
rect 1104 37018 18860 37040
rect 1104 36966 6880 37018
rect 6932 36966 6944 37018
rect 6996 36966 7008 37018
rect 7060 36966 7072 37018
rect 7124 36966 7136 37018
rect 7188 36966 12811 37018
rect 12863 36966 12875 37018
rect 12927 36966 12939 37018
rect 12991 36966 13003 37018
rect 13055 36966 13067 37018
rect 13119 36966 18860 37018
rect 1104 36944 18860 36966
rect 2869 36907 2927 36913
rect 2869 36873 2881 36907
rect 2915 36904 2927 36907
rect 3786 36904 3792 36916
rect 2915 36876 3792 36904
rect 2915 36873 2927 36876
rect 2869 36867 2927 36873
rect 3786 36864 3792 36876
rect 3844 36864 3850 36916
rect 4249 36907 4307 36913
rect 4249 36873 4261 36907
rect 4295 36904 4307 36907
rect 4982 36904 4988 36916
rect 4295 36876 4988 36904
rect 4295 36873 4307 36876
rect 4249 36867 4307 36873
rect 4982 36864 4988 36876
rect 5040 36864 5046 36916
rect 6546 36904 6552 36916
rect 6507 36876 6552 36904
rect 6546 36864 6552 36876
rect 6604 36864 6610 36916
rect 7101 36907 7159 36913
rect 7101 36873 7113 36907
rect 7147 36904 7159 36907
rect 7466 36904 7472 36916
rect 7147 36876 7472 36904
rect 7147 36873 7159 36876
rect 7101 36867 7159 36873
rect 4706 36836 4712 36848
rect 4667 36808 4712 36836
rect 4706 36796 4712 36808
rect 4764 36796 4770 36848
rect 5169 36839 5227 36845
rect 5169 36805 5181 36839
rect 5215 36836 5227 36839
rect 5442 36836 5448 36848
rect 5215 36808 5448 36836
rect 5215 36805 5227 36808
rect 5169 36799 5227 36805
rect 5442 36796 5448 36808
rect 5500 36796 5506 36848
rect 2501 36771 2559 36777
rect 2501 36737 2513 36771
rect 2547 36768 2559 36771
rect 2774 36768 2780 36780
rect 2547 36740 2780 36768
rect 2547 36737 2559 36740
rect 2501 36731 2559 36737
rect 2774 36728 2780 36740
rect 2832 36728 2838 36780
rect 3881 36771 3939 36777
rect 3881 36737 3893 36771
rect 3927 36768 3939 36771
rect 3927 36740 5028 36768
rect 3927 36737 3939 36740
rect 3881 36731 3939 36737
rect 2593 36703 2651 36709
rect 2593 36669 2605 36703
rect 2639 36700 2651 36703
rect 2682 36700 2688 36712
rect 2639 36672 2688 36700
rect 2639 36669 2651 36672
rect 2593 36663 2651 36669
rect 2682 36660 2688 36672
rect 2740 36700 2746 36712
rect 2958 36700 2964 36712
rect 2740 36672 2964 36700
rect 2740 36660 2746 36672
rect 2958 36660 2964 36672
rect 3016 36660 3022 36712
rect 3602 36660 3608 36712
rect 3660 36700 3666 36712
rect 3789 36703 3847 36709
rect 3789 36700 3801 36703
rect 3660 36672 3801 36700
rect 3660 36660 3666 36672
rect 3789 36669 3801 36672
rect 3835 36669 3847 36703
rect 3789 36663 3847 36669
rect 4614 36660 4620 36712
rect 4672 36700 4678 36712
rect 4801 36703 4859 36709
rect 4801 36700 4813 36703
rect 4672 36672 4813 36700
rect 4672 36660 4678 36672
rect 4801 36669 4813 36672
rect 4847 36669 4859 36703
rect 5000 36700 5028 36740
rect 5074 36728 5080 36780
rect 5132 36768 5138 36780
rect 5132 36740 5177 36768
rect 5132 36728 5138 36740
rect 5350 36728 5356 36780
rect 5408 36768 5414 36780
rect 5629 36771 5687 36777
rect 5629 36768 5641 36771
rect 5408 36740 5641 36768
rect 5408 36728 5414 36740
rect 5629 36737 5641 36740
rect 5675 36737 5687 36771
rect 5629 36731 5687 36737
rect 6641 36771 6699 36777
rect 6641 36737 6653 36771
rect 6687 36768 6699 36771
rect 7116 36768 7144 36867
rect 7466 36864 7472 36876
rect 7524 36864 7530 36916
rect 10226 36864 10232 36916
rect 10284 36904 10290 36916
rect 10505 36907 10563 36913
rect 10505 36904 10517 36907
rect 10284 36876 10517 36904
rect 10284 36864 10290 36876
rect 10505 36873 10517 36876
rect 10551 36873 10563 36907
rect 10505 36867 10563 36873
rect 13449 36907 13507 36913
rect 13449 36873 13461 36907
rect 13495 36904 13507 36907
rect 13814 36904 13820 36916
rect 13495 36876 13820 36904
rect 13495 36873 13507 36876
rect 13449 36867 13507 36873
rect 13814 36864 13820 36876
rect 13872 36864 13878 36916
rect 7374 36796 7380 36848
rect 7432 36836 7438 36848
rect 8110 36836 8116 36848
rect 7432 36808 8116 36836
rect 7432 36796 7438 36808
rect 8110 36796 8116 36808
rect 8168 36836 8174 36848
rect 8168 36808 8524 36836
rect 8168 36796 8174 36808
rect 6687 36740 7144 36768
rect 6687 36737 6699 36740
rect 6641 36731 6699 36737
rect 7834 36728 7840 36780
rect 7892 36768 7898 36780
rect 8496 36777 8524 36808
rect 9398 36777 9404 36780
rect 8214 36771 8272 36777
rect 8214 36768 8226 36771
rect 7892 36740 8226 36768
rect 7892 36728 7898 36740
rect 8214 36737 8226 36740
rect 8260 36737 8272 36771
rect 8214 36731 8272 36737
rect 8481 36771 8539 36777
rect 8481 36737 8493 36771
rect 8527 36768 8539 36771
rect 9125 36771 9183 36777
rect 9125 36768 9137 36771
rect 8527 36740 9137 36768
rect 8527 36737 8539 36740
rect 8481 36731 8539 36737
rect 9125 36737 9137 36740
rect 9171 36737 9183 36771
rect 9392 36768 9404 36777
rect 9359 36740 9404 36768
rect 9125 36731 9183 36737
rect 9392 36731 9404 36740
rect 9398 36728 9404 36731
rect 9456 36728 9462 36780
rect 12710 36728 12716 36780
rect 12768 36768 12774 36780
rect 13541 36771 13599 36777
rect 13541 36768 13553 36771
rect 12768 36740 13553 36768
rect 12768 36728 12774 36740
rect 13541 36737 13553 36740
rect 13587 36737 13599 36771
rect 13541 36731 13599 36737
rect 15378 36728 15384 36780
rect 15436 36768 15442 36780
rect 15562 36768 15568 36780
rect 15436 36740 15568 36768
rect 15436 36728 15442 36740
rect 15562 36728 15568 36740
rect 15620 36728 15626 36780
rect 5721 36703 5779 36709
rect 5721 36700 5733 36703
rect 5000 36672 5733 36700
rect 4801 36663 4859 36669
rect 5644 36644 5672 36672
rect 5721 36669 5733 36672
rect 5767 36669 5779 36703
rect 5721 36663 5779 36669
rect 15749 36703 15807 36709
rect 15749 36669 15761 36703
rect 15795 36700 15807 36703
rect 16574 36700 16580 36712
rect 15795 36672 16580 36700
rect 15795 36669 15807 36672
rect 15749 36663 15807 36669
rect 16574 36660 16580 36672
rect 16632 36700 16638 36712
rect 17402 36700 17408 36712
rect 16632 36672 17408 36700
rect 16632 36660 16638 36672
rect 17402 36660 17408 36672
rect 17460 36660 17466 36712
rect 5626 36592 5632 36644
rect 5684 36592 5690 36644
rect 4890 36564 4896 36576
rect 4851 36536 4896 36564
rect 4890 36524 4896 36536
rect 4948 36524 4954 36576
rect 15378 36564 15384 36576
rect 15339 36536 15384 36564
rect 15378 36524 15384 36536
rect 15436 36524 15442 36576
rect 1104 36474 18860 36496
rect 1104 36422 3915 36474
rect 3967 36422 3979 36474
rect 4031 36422 4043 36474
rect 4095 36422 4107 36474
rect 4159 36422 4171 36474
rect 4223 36422 9846 36474
rect 9898 36422 9910 36474
rect 9962 36422 9974 36474
rect 10026 36422 10038 36474
rect 10090 36422 10102 36474
rect 10154 36422 15776 36474
rect 15828 36422 15840 36474
rect 15892 36422 15904 36474
rect 15956 36422 15968 36474
rect 16020 36422 16032 36474
rect 16084 36422 18860 36474
rect 1104 36400 18860 36422
rect 3142 36320 3148 36372
rect 3200 36360 3206 36372
rect 3881 36363 3939 36369
rect 3881 36360 3893 36363
rect 3200 36332 3893 36360
rect 3200 36320 3206 36332
rect 3881 36329 3893 36332
rect 3927 36329 3939 36363
rect 3881 36323 3939 36329
rect 4433 36363 4491 36369
rect 4433 36329 4445 36363
rect 4479 36360 4491 36363
rect 4890 36360 4896 36372
rect 4479 36332 4896 36360
rect 4479 36329 4491 36332
rect 4433 36323 4491 36329
rect 4890 36320 4896 36332
rect 4948 36320 4954 36372
rect 7834 36360 7840 36372
rect 7795 36332 7840 36360
rect 7834 36320 7840 36332
rect 7892 36320 7898 36372
rect 10502 36320 10508 36372
rect 10560 36360 10566 36372
rect 10781 36363 10839 36369
rect 10781 36360 10793 36363
rect 10560 36332 10793 36360
rect 10560 36320 10566 36332
rect 10781 36329 10793 36332
rect 10827 36329 10839 36363
rect 10781 36323 10839 36329
rect 8205 36295 8263 36301
rect 8205 36261 8217 36295
rect 8251 36292 8263 36295
rect 8386 36292 8392 36304
rect 8251 36264 8392 36292
rect 8251 36261 8263 36264
rect 8205 36255 8263 36261
rect 8386 36252 8392 36264
rect 8444 36252 8450 36304
rect 16117 36295 16175 36301
rect 16117 36261 16129 36295
rect 16163 36292 16175 36295
rect 16574 36292 16580 36304
rect 16163 36264 16580 36292
rect 16163 36261 16175 36264
rect 16117 36255 16175 36261
rect 16574 36252 16580 36264
rect 16632 36252 16638 36304
rect 4522 36224 4528 36236
rect 3804 36196 4528 36224
rect 3804 36165 3832 36196
rect 4522 36184 4528 36196
rect 4580 36184 4586 36236
rect 8110 36184 8116 36236
rect 8168 36224 8174 36236
rect 8941 36227 8999 36233
rect 8941 36224 8953 36227
rect 8168 36196 8953 36224
rect 8168 36184 8174 36196
rect 8941 36193 8953 36196
rect 8987 36193 8999 36227
rect 8941 36187 8999 36193
rect 3789 36159 3847 36165
rect 3789 36125 3801 36159
rect 3835 36125 3847 36159
rect 3789 36119 3847 36125
rect 3973 36159 4031 36165
rect 3973 36125 3985 36159
rect 4019 36125 4031 36159
rect 3973 36119 4031 36125
rect 4433 36159 4491 36165
rect 4433 36125 4445 36159
rect 4479 36125 4491 36159
rect 4433 36119 4491 36125
rect 4617 36159 4675 36165
rect 4617 36125 4629 36159
rect 4663 36156 4675 36159
rect 5350 36156 5356 36168
rect 4663 36128 5356 36156
rect 4663 36125 4675 36128
rect 4617 36119 4675 36125
rect 3602 36048 3608 36100
rect 3660 36088 3666 36100
rect 3988 36088 4016 36119
rect 3660 36060 4016 36088
rect 4448 36088 4476 36119
rect 5350 36116 5356 36128
rect 5408 36116 5414 36168
rect 7926 36116 7932 36168
rect 7984 36156 7990 36168
rect 8021 36159 8079 36165
rect 8021 36156 8033 36159
rect 7984 36128 8033 36156
rect 7984 36116 7990 36128
rect 8021 36125 8033 36128
rect 8067 36125 8079 36159
rect 8021 36119 8079 36125
rect 8294 36116 8300 36168
rect 8352 36156 8358 36168
rect 8352 36128 8397 36156
rect 8352 36116 8358 36128
rect 10594 36116 10600 36168
rect 10652 36156 10658 36168
rect 10781 36159 10839 36165
rect 10781 36156 10793 36159
rect 10652 36128 10793 36156
rect 10652 36116 10658 36128
rect 10781 36125 10793 36128
rect 10827 36125 10839 36159
rect 10962 36156 10968 36168
rect 10923 36128 10968 36156
rect 10781 36119 10839 36125
rect 10962 36116 10968 36128
rect 11020 36116 11026 36168
rect 14918 36156 14924 36168
rect 14879 36128 14924 36156
rect 14918 36116 14924 36128
rect 14976 36116 14982 36168
rect 15105 36159 15163 36165
rect 15105 36125 15117 36159
rect 15151 36156 15163 36159
rect 16482 36156 16488 36168
rect 15151 36128 16488 36156
rect 15151 36125 15163 36128
rect 15105 36119 15163 36125
rect 16482 36116 16488 36128
rect 16540 36116 16546 36168
rect 4798 36088 4804 36100
rect 4448 36060 4804 36088
rect 3660 36048 3666 36060
rect 4798 36048 4804 36060
rect 4856 36048 4862 36100
rect 9214 36097 9220 36100
rect 9208 36051 9220 36097
rect 9272 36088 9278 36100
rect 15841 36091 15899 36097
rect 9272 36060 9308 36088
rect 9214 36048 9220 36051
rect 9272 36048 9278 36060
rect 15841 36057 15853 36091
rect 15887 36088 15899 36091
rect 15887 36060 16574 36088
rect 15887 36057 15899 36060
rect 15841 36051 15899 36057
rect 8846 35980 8852 36032
rect 8904 36020 8910 36032
rect 10321 36023 10379 36029
rect 10321 36020 10333 36023
rect 8904 35992 10333 36020
rect 8904 35980 8910 35992
rect 10321 35989 10333 35992
rect 10367 35989 10379 36023
rect 14734 36020 14740 36032
rect 14695 35992 14740 36020
rect 10321 35983 10379 35989
rect 14734 35980 14740 35992
rect 14792 35980 14798 36032
rect 15194 35980 15200 36032
rect 15252 36020 15258 36032
rect 15565 36023 15623 36029
rect 15565 36020 15577 36023
rect 15252 35992 15577 36020
rect 15252 35980 15258 35992
rect 15565 35989 15577 35992
rect 15611 35989 15623 36023
rect 15565 35983 15623 35989
rect 15654 35980 15660 36032
rect 15712 36020 15718 36032
rect 15749 36023 15807 36029
rect 15749 36020 15761 36023
rect 15712 35992 15761 36020
rect 15712 35980 15718 35992
rect 15749 35989 15761 35992
rect 15795 35989 15807 36023
rect 15749 35983 15807 35989
rect 15933 36023 15991 36029
rect 15933 35989 15945 36023
rect 15979 36020 15991 36023
rect 16114 36020 16120 36032
rect 15979 35992 16120 36020
rect 15979 35989 15991 35992
rect 15933 35983 15991 35989
rect 16114 35980 16120 35992
rect 16172 35980 16178 36032
rect 16546 36020 16574 36060
rect 16758 36020 16764 36032
rect 16546 35992 16764 36020
rect 16758 35980 16764 35992
rect 16816 35980 16822 36032
rect 1104 35930 18860 35952
rect 1104 35878 6880 35930
rect 6932 35878 6944 35930
rect 6996 35878 7008 35930
rect 7060 35878 7072 35930
rect 7124 35878 7136 35930
rect 7188 35878 12811 35930
rect 12863 35878 12875 35930
rect 12927 35878 12939 35930
rect 12991 35878 13003 35930
rect 13055 35878 13067 35930
rect 13119 35878 18860 35930
rect 1104 35856 18860 35878
rect 9125 35819 9183 35825
rect 9125 35785 9137 35819
rect 9171 35816 9183 35819
rect 9214 35816 9220 35828
rect 9171 35788 9220 35816
rect 9171 35785 9183 35788
rect 9125 35779 9183 35785
rect 9214 35776 9220 35788
rect 9272 35776 9278 35828
rect 14277 35819 14335 35825
rect 14277 35785 14289 35819
rect 14323 35785 14335 35819
rect 14277 35779 14335 35785
rect 14292 35748 14320 35779
rect 16482 35776 16488 35828
rect 16540 35816 16546 35828
rect 17129 35819 17187 35825
rect 17129 35816 17141 35819
rect 16540 35788 17141 35816
rect 16540 35776 16546 35788
rect 17129 35785 17141 35788
rect 17175 35785 17187 35819
rect 17129 35779 17187 35785
rect 14982 35751 15040 35757
rect 14982 35748 14994 35751
rect 14292 35720 14994 35748
rect 14982 35717 14994 35720
rect 15028 35717 15040 35751
rect 14982 35711 15040 35717
rect 4522 35640 4528 35692
rect 4580 35680 4586 35692
rect 5077 35683 5135 35689
rect 5077 35680 5089 35683
rect 4580 35652 5089 35680
rect 4580 35640 4586 35652
rect 5077 35649 5089 35652
rect 5123 35649 5135 35683
rect 5077 35643 5135 35649
rect 8846 35640 8852 35692
rect 8904 35680 8910 35692
rect 9398 35680 9404 35692
rect 8904 35652 9404 35680
rect 8904 35640 8910 35652
rect 9398 35640 9404 35652
rect 9456 35640 9462 35692
rect 9493 35683 9551 35689
rect 9493 35649 9505 35683
rect 9539 35649 9551 35683
rect 9493 35643 9551 35649
rect 1394 35612 1400 35624
rect 1355 35584 1400 35612
rect 1394 35572 1400 35584
rect 1452 35572 1458 35624
rect 1670 35612 1676 35624
rect 1631 35584 1676 35612
rect 1670 35572 1676 35584
rect 1728 35572 1734 35624
rect 8386 35572 8392 35624
rect 8444 35612 8450 35624
rect 9508 35612 9536 35643
rect 9582 35640 9588 35692
rect 9640 35680 9646 35692
rect 9769 35683 9827 35689
rect 9640 35652 9685 35680
rect 9640 35640 9646 35652
rect 9769 35649 9781 35683
rect 9815 35680 9827 35683
rect 10594 35680 10600 35692
rect 9815 35652 10600 35680
rect 9815 35649 9827 35652
rect 9769 35643 9827 35649
rect 10594 35640 10600 35652
rect 10652 35680 10658 35692
rect 11146 35680 11152 35692
rect 10652 35652 11152 35680
rect 10652 35640 10658 35652
rect 11146 35640 11152 35652
rect 11204 35640 11210 35692
rect 14093 35683 14151 35689
rect 14093 35649 14105 35683
rect 14139 35680 14151 35683
rect 15378 35680 15384 35692
rect 14139 35652 15384 35680
rect 14139 35649 14151 35652
rect 14093 35643 14151 35649
rect 15378 35640 15384 35652
rect 15436 35640 15442 35692
rect 16669 35683 16727 35689
rect 16669 35680 16681 35683
rect 16132 35652 16681 35680
rect 9674 35612 9680 35624
rect 8444 35584 9680 35612
rect 8444 35572 8450 35584
rect 9674 35572 9680 35584
rect 9732 35572 9738 35624
rect 13814 35572 13820 35624
rect 13872 35612 13878 35624
rect 14550 35612 14556 35624
rect 13872 35584 14556 35612
rect 13872 35572 13878 35584
rect 14550 35572 14556 35584
rect 14608 35612 14614 35624
rect 14737 35615 14795 35621
rect 14737 35612 14749 35615
rect 14608 35584 14749 35612
rect 14608 35572 14614 35584
rect 14737 35581 14749 35584
rect 14783 35581 14795 35615
rect 14737 35575 14795 35581
rect 5169 35479 5227 35485
rect 5169 35445 5181 35479
rect 5215 35476 5227 35479
rect 5718 35476 5724 35488
rect 5215 35448 5724 35476
rect 5215 35445 5227 35448
rect 5169 35439 5227 35445
rect 5718 35436 5724 35448
rect 5776 35436 5782 35488
rect 15654 35436 15660 35488
rect 15712 35476 15718 35488
rect 16132 35485 16160 35652
rect 16669 35649 16681 35652
rect 16715 35649 16727 35683
rect 16669 35643 16727 35649
rect 16945 35683 17003 35689
rect 16945 35649 16957 35683
rect 16991 35680 17003 35683
rect 17402 35680 17408 35692
rect 16991 35652 17408 35680
rect 16991 35649 17003 35652
rect 16945 35643 17003 35649
rect 17402 35640 17408 35652
rect 17460 35640 17466 35692
rect 16758 35612 16764 35624
rect 16719 35584 16764 35612
rect 16758 35572 16764 35584
rect 16816 35572 16822 35624
rect 16117 35479 16175 35485
rect 16117 35476 16129 35479
rect 15712 35448 16129 35476
rect 15712 35436 15718 35448
rect 16117 35445 16129 35448
rect 16163 35445 16175 35479
rect 16117 35439 16175 35445
rect 16298 35436 16304 35488
rect 16356 35476 16362 35488
rect 16669 35479 16727 35485
rect 16669 35476 16681 35479
rect 16356 35448 16681 35476
rect 16356 35436 16362 35448
rect 16669 35445 16681 35448
rect 16715 35445 16727 35479
rect 16669 35439 16727 35445
rect 1104 35386 18860 35408
rect 1104 35334 3915 35386
rect 3967 35334 3979 35386
rect 4031 35334 4043 35386
rect 4095 35334 4107 35386
rect 4159 35334 4171 35386
rect 4223 35334 9846 35386
rect 9898 35334 9910 35386
rect 9962 35334 9974 35386
rect 10026 35334 10038 35386
rect 10090 35334 10102 35386
rect 10154 35334 15776 35386
rect 15828 35334 15840 35386
rect 15892 35334 15904 35386
rect 15956 35334 15968 35386
rect 16020 35334 16032 35386
rect 16084 35334 18860 35386
rect 1104 35312 18860 35334
rect 16758 35272 16764 35284
rect 16719 35244 16764 35272
rect 16758 35232 16764 35244
rect 16816 35232 16822 35284
rect 7282 35164 7288 35216
rect 7340 35204 7346 35216
rect 7929 35207 7987 35213
rect 7929 35204 7941 35207
rect 7340 35176 7941 35204
rect 7340 35164 7346 35176
rect 7929 35173 7941 35176
rect 7975 35173 7987 35207
rect 15194 35204 15200 35216
rect 7929 35167 7987 35173
rect 14476 35176 15200 35204
rect 14366 35068 14372 35080
rect 14327 35040 14372 35068
rect 14366 35028 14372 35040
rect 14424 35028 14430 35080
rect 14476 35077 14504 35176
rect 15194 35164 15200 35176
rect 15252 35164 15258 35216
rect 14550 35096 14556 35148
rect 14608 35136 14614 35148
rect 15381 35139 15439 35145
rect 15381 35136 15393 35139
rect 14608 35108 15393 35136
rect 14608 35096 14614 35108
rect 15381 35105 15393 35108
rect 15427 35105 15439 35139
rect 15381 35099 15439 35105
rect 14734 35077 14740 35080
rect 14461 35071 14519 35077
rect 14461 35037 14473 35071
rect 14507 35037 14519 35071
rect 14461 35031 14519 35037
rect 14691 35071 14740 35077
rect 14691 35037 14703 35071
rect 14737 35037 14740 35071
rect 14691 35031 14740 35037
rect 14734 35028 14740 35031
rect 14792 35028 14798 35080
rect 14826 35028 14832 35080
rect 14884 35068 14890 35080
rect 14884 35040 14929 35068
rect 14884 35028 14890 35040
rect 8113 35003 8171 35009
rect 8113 34969 8125 35003
rect 8159 35000 8171 35003
rect 10410 35000 10416 35012
rect 8159 34972 10416 35000
rect 8159 34969 8171 34972
rect 8113 34963 8171 34969
rect 10410 34960 10416 34972
rect 10468 34960 10474 35012
rect 14553 35003 14611 35009
rect 14553 34969 14565 35003
rect 14599 34969 14611 35003
rect 14553 34963 14611 34969
rect 15648 35003 15706 35009
rect 15648 34969 15660 35003
rect 15694 35000 15706 35003
rect 16666 35000 16672 35012
rect 15694 34972 16672 35000
rect 15694 34969 15706 34972
rect 15648 34963 15706 34969
rect 14182 34932 14188 34944
rect 14143 34904 14188 34932
rect 14182 34892 14188 34904
rect 14240 34892 14246 34944
rect 14568 34932 14596 34963
rect 16666 34960 16672 34972
rect 16724 34960 16730 35012
rect 16298 34932 16304 34944
rect 14568 34904 16304 34932
rect 16298 34892 16304 34904
rect 16356 34892 16362 34944
rect 1104 34842 18860 34864
rect 1104 34790 6880 34842
rect 6932 34790 6944 34842
rect 6996 34790 7008 34842
rect 7060 34790 7072 34842
rect 7124 34790 7136 34842
rect 7188 34790 12811 34842
rect 12863 34790 12875 34842
rect 12927 34790 12939 34842
rect 12991 34790 13003 34842
rect 13055 34790 13067 34842
rect 13119 34790 18860 34842
rect 1104 34768 18860 34790
rect 10410 34728 10416 34740
rect 10371 34700 10416 34728
rect 10410 34688 10416 34700
rect 10468 34728 10474 34740
rect 16666 34728 16672 34740
rect 10468 34700 12572 34728
rect 16627 34700 16672 34728
rect 10468 34688 10474 34700
rect 12544 34669 12572 34700
rect 16666 34688 16672 34700
rect 16724 34688 16730 34740
rect 12529 34663 12587 34669
rect 12529 34629 12541 34663
rect 12575 34629 12587 34663
rect 12529 34623 12587 34629
rect 14182 34620 14188 34672
rect 14240 34660 14246 34672
rect 14286 34663 14344 34669
rect 14286 34660 14298 34663
rect 14240 34632 14298 34660
rect 14240 34620 14246 34632
rect 14286 34629 14298 34632
rect 14332 34629 14344 34663
rect 14286 34623 14344 34629
rect 10502 34592 10508 34604
rect 10463 34564 10508 34592
rect 10502 34552 10508 34564
rect 10560 34552 10566 34604
rect 11790 34592 11796 34604
rect 11751 34564 11796 34592
rect 11790 34552 11796 34564
rect 11848 34552 11854 34604
rect 11977 34595 12035 34601
rect 11977 34561 11989 34595
rect 12023 34561 12035 34595
rect 14550 34592 14556 34604
rect 14511 34564 14556 34592
rect 11977 34555 12035 34561
rect 11514 34484 11520 34536
rect 11572 34524 11578 34536
rect 11992 34524 12020 34555
rect 14550 34552 14556 34564
rect 14608 34552 14614 34604
rect 15289 34595 15347 34601
rect 15289 34561 15301 34595
rect 15335 34592 15347 34595
rect 15562 34592 15568 34604
rect 15335 34564 15568 34592
rect 15335 34561 15347 34564
rect 15289 34555 15347 34561
rect 15562 34552 15568 34564
rect 15620 34552 15626 34604
rect 16850 34592 16856 34604
rect 16811 34564 16856 34592
rect 16850 34552 16856 34564
rect 16908 34552 16914 34604
rect 12710 34524 12716 34536
rect 11572 34496 12020 34524
rect 12671 34496 12716 34524
rect 11572 34484 11578 34496
rect 12710 34484 12716 34496
rect 12768 34484 12774 34536
rect 15010 34524 15016 34536
rect 14971 34496 15016 34524
rect 15010 34484 15016 34496
rect 15068 34484 15074 34536
rect 11974 34388 11980 34400
rect 11935 34360 11980 34388
rect 11974 34348 11980 34360
rect 12032 34348 12038 34400
rect 13170 34388 13176 34400
rect 13131 34360 13176 34388
rect 13170 34348 13176 34360
rect 13228 34348 13234 34400
rect 1104 34298 18860 34320
rect 1104 34246 3915 34298
rect 3967 34246 3979 34298
rect 4031 34246 4043 34298
rect 4095 34246 4107 34298
rect 4159 34246 4171 34298
rect 4223 34246 9846 34298
rect 9898 34246 9910 34298
rect 9962 34246 9974 34298
rect 10026 34246 10038 34298
rect 10090 34246 10102 34298
rect 10154 34246 15776 34298
rect 15828 34246 15840 34298
rect 15892 34246 15904 34298
rect 15956 34246 15968 34298
rect 16020 34246 16032 34298
rect 16084 34246 18860 34298
rect 1104 34224 18860 34246
rect 7837 34187 7895 34193
rect 7837 34153 7849 34187
rect 7883 34184 7895 34187
rect 8018 34184 8024 34196
rect 7883 34156 8024 34184
rect 7883 34153 7895 34156
rect 7837 34147 7895 34153
rect 8018 34144 8024 34156
rect 8076 34144 8082 34196
rect 14277 34187 14335 34193
rect 14277 34153 14289 34187
rect 14323 34184 14335 34187
rect 14826 34184 14832 34196
rect 14323 34156 14832 34184
rect 14323 34153 14335 34156
rect 14277 34147 14335 34153
rect 5902 33940 5908 33992
rect 5960 33980 5966 33992
rect 5997 33983 6055 33989
rect 5997 33980 6009 33983
rect 5960 33952 6009 33980
rect 5960 33940 5966 33952
rect 5997 33949 6009 33952
rect 6043 33949 6055 33983
rect 5997 33943 6055 33949
rect 6089 33983 6147 33989
rect 6089 33949 6101 33983
rect 6135 33980 6147 33983
rect 6454 33980 6460 33992
rect 6135 33952 6460 33980
rect 6135 33949 6147 33952
rect 6089 33943 6147 33949
rect 6454 33940 6460 33952
rect 6512 33980 6518 33992
rect 6549 33983 6607 33989
rect 6549 33980 6561 33983
rect 6512 33952 6561 33980
rect 6512 33940 6518 33952
rect 6549 33949 6561 33952
rect 6595 33949 6607 33983
rect 6549 33943 6607 33949
rect 6733 33983 6791 33989
rect 6733 33949 6745 33983
rect 6779 33980 6791 33983
rect 7558 33980 7564 33992
rect 6779 33952 7564 33980
rect 6779 33949 6791 33952
rect 6733 33943 6791 33949
rect 7558 33940 7564 33952
rect 7616 33940 7622 33992
rect 7929 33983 7987 33989
rect 7929 33949 7941 33983
rect 7975 33980 7987 33983
rect 9122 33980 9128 33992
rect 7975 33952 9128 33980
rect 7975 33949 7987 33952
rect 7929 33943 7987 33949
rect 9122 33940 9128 33952
rect 9180 33940 9186 33992
rect 13354 33980 13360 33992
rect 13315 33952 13360 33980
rect 13354 33940 13360 33952
rect 13412 33940 13418 33992
rect 14090 33980 14096 33992
rect 14051 33952 14096 33980
rect 14090 33940 14096 33952
rect 14148 33940 14154 33992
rect 5813 33915 5871 33921
rect 5813 33881 5825 33915
rect 5859 33912 5871 33915
rect 7466 33912 7472 33924
rect 5859 33884 7472 33912
rect 5859 33881 5871 33884
rect 5813 33875 5871 33881
rect 7466 33872 7472 33884
rect 7524 33912 7530 33924
rect 8018 33912 8024 33924
rect 7524 33884 8024 33912
rect 7524 33872 7530 33884
rect 8018 33872 8024 33884
rect 8076 33872 8082 33924
rect 13112 33915 13170 33921
rect 13112 33881 13124 33915
rect 13158 33912 13170 33915
rect 14292 33912 14320 34147
rect 14826 34144 14832 34156
rect 14884 34144 14890 34196
rect 16025 34187 16083 34193
rect 16025 34153 16037 34187
rect 16071 34184 16083 34187
rect 16850 34184 16856 34196
rect 16071 34156 16856 34184
rect 16071 34153 16083 34156
rect 16025 34147 16083 34153
rect 16850 34144 16856 34156
rect 16908 34144 16914 34196
rect 15654 34048 15660 34060
rect 15615 34020 15660 34048
rect 15654 34008 15660 34020
rect 15712 34008 15718 34060
rect 15841 33983 15899 33989
rect 15841 33949 15853 33983
rect 15887 33949 15899 33983
rect 15841 33943 15899 33949
rect 13158 33884 14320 33912
rect 13158 33881 13170 33884
rect 13112 33875 13170 33881
rect 15378 33872 15384 33924
rect 15436 33912 15442 33924
rect 15856 33912 15884 33943
rect 15436 33884 15884 33912
rect 15436 33872 15442 33884
rect 5902 33844 5908 33856
rect 5960 33853 5966 33856
rect 5869 33816 5908 33844
rect 5902 33804 5908 33816
rect 5960 33807 5969 33853
rect 6638 33844 6644 33856
rect 6599 33816 6644 33844
rect 5960 33804 5966 33807
rect 6638 33804 6644 33816
rect 6696 33804 6702 33856
rect 11790 33804 11796 33856
rect 11848 33844 11854 33856
rect 11977 33847 12035 33853
rect 11977 33844 11989 33847
rect 11848 33816 11989 33844
rect 11848 33804 11854 33816
rect 11977 33813 11989 33816
rect 12023 33813 12035 33847
rect 11977 33807 12035 33813
rect 1104 33754 18860 33776
rect 1104 33702 6880 33754
rect 6932 33702 6944 33754
rect 6996 33702 7008 33754
rect 7060 33702 7072 33754
rect 7124 33702 7136 33754
rect 7188 33702 12811 33754
rect 12863 33702 12875 33754
rect 12927 33702 12939 33754
rect 12991 33702 13003 33754
rect 13055 33702 13067 33754
rect 13119 33702 18860 33754
rect 1104 33680 18860 33702
rect 10965 33643 11023 33649
rect 10965 33609 10977 33643
rect 11011 33640 11023 33643
rect 11011 33612 12296 33640
rect 11011 33609 11023 33612
rect 10965 33603 11023 33609
rect 5902 33532 5908 33584
rect 5960 33572 5966 33584
rect 5960 33544 6592 33572
rect 5960 33532 5966 33544
rect 6564 33513 6592 33544
rect 7282 33532 7288 33584
rect 7340 33572 7346 33584
rect 7561 33575 7619 33581
rect 7561 33572 7573 33575
rect 7340 33544 7573 33572
rect 7340 33532 7346 33544
rect 7561 33541 7573 33544
rect 7607 33541 7619 33575
rect 7561 33535 7619 33541
rect 8294 33532 8300 33584
rect 8352 33572 8358 33584
rect 8389 33575 8447 33581
rect 8389 33572 8401 33575
rect 8352 33544 8401 33572
rect 8352 33532 8358 33544
rect 8389 33541 8401 33544
rect 8435 33541 8447 33575
rect 11790 33572 11796 33584
rect 8389 33535 8447 33541
rect 10704 33544 11796 33572
rect 4700 33507 4758 33513
rect 4700 33473 4712 33507
rect 4746 33504 4758 33507
rect 6365 33507 6423 33513
rect 6365 33504 6377 33507
rect 4746 33476 6377 33504
rect 4746 33473 4758 33476
rect 4700 33467 4758 33473
rect 6365 33473 6377 33476
rect 6411 33473 6423 33507
rect 6365 33467 6423 33473
rect 6549 33507 6607 33513
rect 6549 33473 6561 33507
rect 6595 33473 6607 33507
rect 8110 33504 8116 33516
rect 8071 33476 8116 33504
rect 6549 33467 6607 33473
rect 8110 33464 8116 33476
rect 8168 33464 8174 33516
rect 8202 33464 8208 33516
rect 8260 33504 8266 33516
rect 10704 33513 10732 33544
rect 11790 33532 11796 33544
rect 11848 33532 11854 33584
rect 12268 33516 12296 33612
rect 13170 33572 13176 33584
rect 13131 33544 13176 33572
rect 13170 33532 13176 33544
rect 13228 33532 13234 33584
rect 8849 33507 8907 33513
rect 8260 33476 8305 33504
rect 8260 33464 8266 33476
rect 8849 33473 8861 33507
rect 8895 33473 8907 33507
rect 8849 33467 8907 33473
rect 10689 33507 10747 33513
rect 10689 33473 10701 33507
rect 10735 33473 10747 33507
rect 10689 33467 10747 33473
rect 10781 33507 10839 33513
rect 10781 33473 10793 33507
rect 10827 33504 10839 33507
rect 11514 33504 11520 33516
rect 10827 33476 11520 33504
rect 10827 33473 10839 33476
rect 10781 33467 10839 33473
rect 4433 33439 4491 33445
rect 4433 33405 4445 33439
rect 4479 33405 4491 33439
rect 4433 33399 4491 33405
rect 4448 33312 4476 33399
rect 5810 33396 5816 33448
rect 5868 33436 5874 33448
rect 6825 33439 6883 33445
rect 6825 33436 6837 33439
rect 5868 33408 6837 33436
rect 5868 33396 5874 33408
rect 6825 33405 6837 33408
rect 6871 33405 6883 33439
rect 8864 33436 8892 33467
rect 11514 33464 11520 33476
rect 11572 33464 11578 33516
rect 11885 33507 11943 33513
rect 11885 33473 11897 33507
rect 11931 33473 11943 33507
rect 11885 33467 11943 33473
rect 6825 33399 6883 33405
rect 8404 33408 8892 33436
rect 9125 33439 9183 33445
rect 7374 33368 7380 33380
rect 5368 33340 7380 33368
rect 4430 33300 4436 33312
rect 4343 33272 4436 33300
rect 4430 33260 4436 33272
rect 4488 33300 4494 33312
rect 5368 33300 5396 33340
rect 7374 33328 7380 33340
rect 7432 33328 7438 33380
rect 8404 33377 8432 33408
rect 9125 33405 9137 33439
rect 9171 33436 9183 33439
rect 9214 33436 9220 33448
rect 9171 33408 9220 33436
rect 9171 33405 9183 33408
rect 9125 33399 9183 33405
rect 9214 33396 9220 33408
rect 9272 33436 9278 33448
rect 10410 33436 10416 33448
rect 9272 33408 10416 33436
rect 9272 33396 9278 33408
rect 10410 33396 10416 33408
rect 10468 33396 10474 33448
rect 11900 33436 11928 33467
rect 11974 33464 11980 33516
rect 12032 33504 12038 33516
rect 12032 33476 12077 33504
rect 12032 33464 12038 33476
rect 12250 33464 12256 33516
rect 12308 33504 12314 33516
rect 12308 33476 12401 33504
rect 12308 33464 12314 33476
rect 13998 33464 14004 33516
rect 14056 33504 14062 33516
rect 14366 33504 14372 33516
rect 14056 33476 14372 33504
rect 14056 33464 14062 33476
rect 14366 33464 14372 33476
rect 14424 33504 14430 33516
rect 14737 33507 14795 33513
rect 14737 33504 14749 33507
rect 14424 33476 14749 33504
rect 14424 33464 14430 33476
rect 14737 33473 14749 33476
rect 14783 33473 14795 33507
rect 14737 33467 14795 33473
rect 12066 33436 12072 33448
rect 11900 33408 12072 33436
rect 12066 33396 12072 33408
rect 12124 33436 12130 33448
rect 12713 33439 12771 33445
rect 12713 33436 12725 33439
rect 12124 33408 12725 33436
rect 12124 33396 12130 33408
rect 12713 33405 12725 33408
rect 12759 33405 12771 33439
rect 15010 33436 15016 33448
rect 14971 33408 15016 33436
rect 12713 33399 12771 33405
rect 15010 33396 15016 33408
rect 15068 33396 15074 33448
rect 8389 33371 8447 33377
rect 8389 33337 8401 33371
rect 8435 33337 8447 33371
rect 8389 33331 8447 33337
rect 8754 33328 8760 33380
rect 8812 33368 8818 33380
rect 9033 33371 9091 33377
rect 9033 33368 9045 33371
rect 8812 33340 9045 33368
rect 8812 33328 8818 33340
rect 9033 33337 9045 33340
rect 9079 33337 9091 33371
rect 9033 33331 9091 33337
rect 12434 33328 12440 33380
rect 12492 33368 12498 33380
rect 12805 33371 12863 33377
rect 12805 33368 12817 33371
rect 12492 33340 12817 33368
rect 12492 33328 12498 33340
rect 12805 33337 12817 33340
rect 12851 33337 12863 33371
rect 12805 33331 12863 33337
rect 5810 33300 5816 33312
rect 4488 33272 5396 33300
rect 5771 33272 5816 33300
rect 4488 33260 4494 33272
rect 5810 33260 5816 33272
rect 5868 33260 5874 33312
rect 6454 33260 6460 33312
rect 6512 33300 6518 33312
rect 6733 33303 6791 33309
rect 6733 33300 6745 33303
rect 6512 33272 6745 33300
rect 6512 33260 6518 33272
rect 6733 33269 6745 33272
rect 6779 33269 6791 33303
rect 8938 33300 8944 33312
rect 8899 33272 8944 33300
rect 6733 33263 6791 33269
rect 8938 33260 8944 33272
rect 8996 33260 9002 33312
rect 10226 33260 10232 33312
rect 10284 33300 10290 33312
rect 11701 33303 11759 33309
rect 11701 33300 11713 33303
rect 10284 33272 11713 33300
rect 10284 33260 10290 33272
rect 11701 33269 11713 33272
rect 11747 33269 11759 33303
rect 11701 33263 11759 33269
rect 11882 33260 11888 33312
rect 11940 33300 11946 33312
rect 12161 33303 12219 33309
rect 12161 33300 12173 33303
rect 11940 33272 12173 33300
rect 11940 33260 11946 33272
rect 12161 33269 12173 33272
rect 12207 33269 12219 33303
rect 12161 33263 12219 33269
rect 1104 33210 18860 33232
rect 1104 33158 3915 33210
rect 3967 33158 3979 33210
rect 4031 33158 4043 33210
rect 4095 33158 4107 33210
rect 4159 33158 4171 33210
rect 4223 33158 9846 33210
rect 9898 33158 9910 33210
rect 9962 33158 9974 33210
rect 10026 33158 10038 33210
rect 10090 33158 10102 33210
rect 10154 33158 15776 33210
rect 15828 33158 15840 33210
rect 15892 33158 15904 33210
rect 15956 33158 15968 33210
rect 16020 33158 16032 33210
rect 16084 33158 18860 33210
rect 1104 33136 18860 33158
rect 4706 33056 4712 33108
rect 4764 33096 4770 33108
rect 8205 33099 8263 33105
rect 4764 33068 6960 33096
rect 4764 33056 4770 33068
rect 5074 33028 5080 33040
rect 3804 33000 5080 33028
rect 3694 32852 3700 32904
rect 3752 32892 3758 32904
rect 3804 32892 3832 33000
rect 5074 32988 5080 33000
rect 5132 32988 5138 33040
rect 6932 33028 6960 33068
rect 8205 33065 8217 33099
rect 8251 33096 8263 33099
rect 8294 33096 8300 33108
rect 8251 33068 8300 33096
rect 8251 33065 8263 33068
rect 8205 33059 8263 33065
rect 8294 33056 8300 33068
rect 8352 33056 8358 33108
rect 8389 33099 8447 33105
rect 8389 33065 8401 33099
rect 8435 33096 8447 33099
rect 8938 33096 8944 33108
rect 8435 33068 8944 33096
rect 8435 33065 8447 33068
rect 8389 33059 8447 33065
rect 8938 33056 8944 33068
rect 8996 33056 9002 33108
rect 10686 33096 10692 33108
rect 9048 33068 10692 33096
rect 9048 33028 9076 33068
rect 10686 33056 10692 33068
rect 10744 33056 10750 33108
rect 11514 33096 11520 33108
rect 11475 33068 11520 33096
rect 11514 33056 11520 33068
rect 11572 33056 11578 33108
rect 14090 33096 14096 33108
rect 14051 33068 14096 33096
rect 14090 33056 14096 33068
rect 14148 33056 14154 33108
rect 6932 33000 9076 33028
rect 9674 32988 9680 33040
rect 9732 33028 9738 33040
rect 10045 33031 10103 33037
rect 10045 33028 10057 33031
rect 9732 33000 10057 33028
rect 9732 32988 9738 33000
rect 10045 32997 10057 33000
rect 10091 32997 10103 33031
rect 10045 32991 10103 32997
rect 10410 32988 10416 33040
rect 10468 33028 10474 33040
rect 10781 33031 10839 33037
rect 10781 33028 10793 33031
rect 10468 33000 10793 33028
rect 10468 32988 10474 33000
rect 10781 32997 10793 33000
rect 10827 32997 10839 33031
rect 10781 32991 10839 32997
rect 3881 32963 3939 32969
rect 3881 32929 3893 32963
rect 3927 32960 3939 32963
rect 4614 32960 4620 32972
rect 3927 32932 4620 32960
rect 3927 32929 3939 32932
rect 3881 32923 3939 32929
rect 4614 32920 4620 32932
rect 4672 32960 4678 32972
rect 5626 32960 5632 32972
rect 4672 32932 4936 32960
rect 4672 32920 4678 32932
rect 3973 32895 4031 32901
rect 3752 32864 3924 32892
rect 3752 32852 3758 32864
rect 3789 32827 3847 32833
rect 3789 32793 3801 32827
rect 3835 32793 3847 32827
rect 3896 32824 3924 32864
rect 3973 32861 3985 32895
rect 4019 32892 4031 32895
rect 4522 32892 4528 32904
rect 4019 32864 4528 32892
rect 4019 32861 4031 32864
rect 3973 32855 4031 32861
rect 4522 32852 4528 32864
rect 4580 32852 4586 32904
rect 4706 32892 4712 32904
rect 4667 32864 4712 32892
rect 4706 32852 4712 32864
rect 4764 32852 4770 32904
rect 4246 32824 4252 32836
rect 3896 32796 4016 32824
rect 4207 32796 4252 32824
rect 3789 32787 3847 32793
rect 3804 32756 3832 32787
rect 3878 32756 3884 32768
rect 3804 32728 3884 32756
rect 3878 32716 3884 32728
rect 3936 32716 3942 32768
rect 3988 32756 4016 32796
rect 4246 32784 4252 32796
rect 4304 32784 4310 32836
rect 4908 32824 4936 32932
rect 5276 32932 5632 32960
rect 4985 32895 5043 32901
rect 4985 32861 4997 32895
rect 5031 32892 5043 32895
rect 5074 32892 5080 32904
rect 5031 32864 5080 32892
rect 5031 32861 5043 32864
rect 4985 32855 5043 32861
rect 5074 32852 5080 32864
rect 5132 32852 5138 32904
rect 5276 32901 5304 32932
rect 5626 32920 5632 32932
rect 5684 32920 5690 32972
rect 8202 32920 8208 32972
rect 8260 32960 8266 32972
rect 9030 32960 9036 32972
rect 8260 32932 9036 32960
rect 8260 32920 8266 32932
rect 9030 32920 9036 32932
rect 9088 32920 9094 32972
rect 10226 32960 10232 32972
rect 9324 32932 10232 32960
rect 5261 32895 5319 32901
rect 5261 32861 5273 32895
rect 5307 32861 5319 32895
rect 5261 32855 5319 32861
rect 5537 32895 5595 32901
rect 5537 32861 5549 32895
rect 5583 32892 5595 32895
rect 5810 32892 5816 32904
rect 5583 32864 5816 32892
rect 5583 32861 5595 32864
rect 5537 32855 5595 32861
rect 5810 32852 5816 32864
rect 5868 32852 5874 32904
rect 5997 32895 6055 32901
rect 5997 32861 6009 32895
rect 6043 32892 6055 32895
rect 7374 32892 7380 32904
rect 6043 32864 7380 32892
rect 6043 32861 6055 32864
rect 5997 32855 6055 32861
rect 7374 32852 7380 32864
rect 7432 32852 7438 32904
rect 8386 32892 8392 32904
rect 8036 32864 8392 32892
rect 6264 32827 6322 32833
rect 4908 32796 6224 32824
rect 6196 32768 6224 32796
rect 6264 32793 6276 32827
rect 6310 32824 6322 32827
rect 6638 32824 6644 32836
rect 6310 32796 6644 32824
rect 6310 32793 6322 32796
rect 6264 32787 6322 32793
rect 6638 32784 6644 32796
rect 6696 32784 6702 32836
rect 8036 32833 8064 32864
rect 8386 32852 8392 32864
rect 8444 32852 8450 32904
rect 9122 32892 9128 32904
rect 9083 32864 9128 32892
rect 9122 32852 9128 32864
rect 9180 32852 9186 32904
rect 9324 32901 9352 32932
rect 10226 32920 10232 32932
rect 10284 32920 10290 32972
rect 13170 32920 13176 32972
rect 13228 32960 13234 32972
rect 14461 32963 14519 32969
rect 14461 32960 14473 32963
rect 13228 32932 14473 32960
rect 13228 32920 13234 32932
rect 14461 32929 14473 32932
rect 14507 32929 14519 32963
rect 15378 32960 15384 32972
rect 15339 32932 15384 32960
rect 14461 32923 14519 32929
rect 15378 32920 15384 32932
rect 15436 32960 15442 32972
rect 16758 32960 16764 32972
rect 15436 32932 16764 32960
rect 15436 32920 15442 32932
rect 16758 32920 16764 32932
rect 16816 32920 16822 32972
rect 9309 32895 9367 32901
rect 9309 32861 9321 32895
rect 9355 32861 9367 32895
rect 9309 32855 9367 32861
rect 12897 32895 12955 32901
rect 12897 32861 12909 32895
rect 12943 32892 12955 32895
rect 13354 32892 13360 32904
rect 12943 32864 13360 32892
rect 12943 32861 12955 32864
rect 12897 32855 12955 32861
rect 13354 32852 13360 32864
rect 13412 32892 13418 32904
rect 13722 32892 13728 32904
rect 13412 32864 13728 32892
rect 13412 32852 13418 32864
rect 13722 32852 13728 32864
rect 13780 32852 13786 32904
rect 14182 32852 14188 32904
rect 14240 32892 14246 32904
rect 14277 32895 14335 32901
rect 14277 32892 14289 32895
rect 14240 32864 14289 32892
rect 14240 32852 14246 32864
rect 14277 32861 14289 32864
rect 14323 32861 14335 32895
rect 14277 32855 14335 32861
rect 15010 32852 15016 32904
rect 15068 32892 15074 32904
rect 15105 32895 15163 32901
rect 15105 32892 15117 32895
rect 15068 32864 15117 32892
rect 15068 32852 15074 32864
rect 15105 32861 15117 32864
rect 15151 32861 15163 32895
rect 15105 32855 15163 32861
rect 8021 32827 8079 32833
rect 8021 32793 8033 32827
rect 8067 32793 8079 32827
rect 8021 32787 8079 32793
rect 8110 32784 8116 32836
rect 8168 32824 8174 32836
rect 8221 32827 8279 32833
rect 8221 32824 8233 32827
rect 8168 32796 8233 32824
rect 8168 32784 8174 32796
rect 8221 32793 8233 32796
rect 8267 32824 8279 32827
rect 8941 32827 8999 32833
rect 8941 32824 8953 32827
rect 8267 32796 8953 32824
rect 8267 32793 8279 32796
rect 8221 32787 8279 32793
rect 8941 32793 8953 32796
rect 8987 32793 8999 32827
rect 8941 32787 8999 32793
rect 10229 32827 10287 32833
rect 10229 32793 10241 32827
rect 10275 32824 10287 32827
rect 10778 32824 10784 32836
rect 10275 32796 10784 32824
rect 10275 32793 10287 32796
rect 10229 32787 10287 32793
rect 10778 32784 10784 32796
rect 10836 32824 10842 32836
rect 10965 32827 11023 32833
rect 10965 32824 10977 32827
rect 10836 32796 10977 32824
rect 10836 32784 10842 32796
rect 10965 32793 10977 32796
rect 11011 32793 11023 32827
rect 12618 32824 12624 32836
rect 12676 32833 12682 32836
rect 12588 32796 12624 32824
rect 10965 32787 11023 32793
rect 12618 32784 12624 32796
rect 12676 32787 12688 32833
rect 12676 32784 12682 32787
rect 4157 32759 4215 32765
rect 4157 32756 4169 32759
rect 3988 32728 4169 32756
rect 4157 32725 4169 32728
rect 4203 32725 4215 32759
rect 4157 32719 4215 32725
rect 4614 32716 4620 32768
rect 4672 32756 4678 32768
rect 4801 32759 4859 32765
rect 4801 32756 4813 32759
rect 4672 32728 4813 32756
rect 4672 32716 4678 32728
rect 4801 32725 4813 32728
rect 4847 32725 4859 32759
rect 4801 32719 4859 32725
rect 6178 32716 6184 32768
rect 6236 32716 6242 32768
rect 7282 32716 7288 32768
rect 7340 32756 7346 32768
rect 7377 32759 7435 32765
rect 7377 32756 7389 32759
rect 7340 32728 7389 32756
rect 7340 32716 7346 32728
rect 7377 32725 7389 32728
rect 7423 32725 7435 32759
rect 7377 32719 7435 32725
rect 1104 32666 18860 32688
rect 1104 32614 6880 32666
rect 6932 32614 6944 32666
rect 6996 32614 7008 32666
rect 7060 32614 7072 32666
rect 7124 32614 7136 32666
rect 7188 32614 12811 32666
rect 12863 32614 12875 32666
rect 12927 32614 12939 32666
rect 12991 32614 13003 32666
rect 13055 32614 13067 32666
rect 13119 32614 18860 32666
rect 1104 32592 18860 32614
rect 6454 32552 6460 32564
rect 6415 32524 6460 32552
rect 6454 32512 6460 32524
rect 6512 32512 6518 32564
rect 6625 32555 6683 32561
rect 6625 32521 6637 32555
rect 6671 32552 6683 32555
rect 7558 32552 7564 32564
rect 6671 32524 7420 32552
rect 7519 32524 7564 32552
rect 6671 32521 6683 32524
rect 6625 32515 6683 32521
rect 4430 32484 4436 32496
rect 3620 32456 4436 32484
rect 3620 32425 3648 32456
rect 4430 32444 4436 32456
rect 4488 32444 4494 32496
rect 5994 32484 6000 32496
rect 5644 32456 6000 32484
rect 3878 32425 3884 32428
rect 3605 32419 3663 32425
rect 3605 32385 3617 32419
rect 3651 32385 3663 32419
rect 3872 32416 3884 32425
rect 3839 32388 3884 32416
rect 3605 32379 3663 32385
rect 3872 32379 3884 32388
rect 3878 32376 3884 32379
rect 3936 32376 3942 32428
rect 5644 32425 5672 32456
rect 5994 32444 6000 32456
rect 6052 32444 6058 32496
rect 6086 32444 6092 32496
rect 6144 32484 6150 32496
rect 6825 32487 6883 32493
rect 6825 32484 6837 32487
rect 6144 32456 6837 32484
rect 6144 32444 6150 32456
rect 6825 32453 6837 32456
rect 6871 32484 6883 32487
rect 7098 32484 7104 32496
rect 6871 32456 7104 32484
rect 6871 32453 6883 32456
rect 6825 32447 6883 32453
rect 7098 32444 7104 32456
rect 7156 32484 7162 32496
rect 7392 32484 7420 32524
rect 7558 32512 7564 32524
rect 7616 32512 7622 32564
rect 8846 32552 8852 32564
rect 8807 32524 8852 32552
rect 8846 32512 8852 32524
rect 8904 32512 8910 32564
rect 10137 32555 10195 32561
rect 10137 32521 10149 32555
rect 10183 32552 10195 32555
rect 10318 32552 10324 32564
rect 10183 32524 10324 32552
rect 10183 32521 10195 32524
rect 10137 32515 10195 32521
rect 10318 32512 10324 32524
rect 10376 32512 10382 32564
rect 11882 32512 11888 32564
rect 11940 32552 11946 32564
rect 13173 32555 13231 32561
rect 13173 32552 13185 32555
rect 11940 32524 13185 32552
rect 11940 32512 11946 32524
rect 13173 32521 13185 32524
rect 13219 32521 13231 32555
rect 13173 32515 13231 32521
rect 7926 32484 7932 32496
rect 7156 32456 7236 32484
rect 7392 32456 7932 32484
rect 7156 32444 7162 32456
rect 5629 32419 5687 32425
rect 5629 32385 5641 32419
rect 5675 32385 5687 32419
rect 5629 32379 5687 32385
rect 5813 32419 5871 32425
rect 5813 32385 5825 32419
rect 5859 32385 5871 32419
rect 7208 32416 7236 32456
rect 7926 32444 7932 32456
rect 7984 32444 7990 32496
rect 8386 32444 8392 32496
rect 8444 32484 8450 32496
rect 8444 32456 8892 32484
rect 8444 32444 8450 32456
rect 7282 32416 7288 32428
rect 7195 32388 7288 32416
rect 5813 32379 5871 32385
rect 5828 32348 5856 32379
rect 7282 32376 7288 32388
rect 7340 32376 7346 32428
rect 8110 32376 8116 32428
rect 8168 32416 8174 32428
rect 8864 32425 8892 32456
rect 9674 32444 9680 32496
rect 9732 32484 9738 32496
rect 10045 32487 10103 32493
rect 10045 32484 10057 32487
rect 9732 32456 10057 32484
rect 9732 32444 9738 32456
rect 10045 32453 10057 32456
rect 10091 32484 10103 32487
rect 10226 32484 10232 32496
rect 10091 32456 10232 32484
rect 10091 32453 10103 32456
rect 10045 32447 10103 32453
rect 10226 32444 10232 32456
rect 10284 32444 10290 32496
rect 10778 32484 10784 32496
rect 10739 32456 10784 32484
rect 10778 32444 10784 32456
rect 10836 32484 10842 32496
rect 11701 32487 11759 32493
rect 11701 32484 11713 32487
rect 10836 32456 11713 32484
rect 10836 32444 10842 32456
rect 11701 32453 11713 32456
rect 11747 32453 11759 32487
rect 11701 32447 11759 32453
rect 12710 32444 12716 32496
rect 12768 32484 12774 32496
rect 13725 32487 13783 32493
rect 13725 32484 13737 32487
rect 12768 32456 13737 32484
rect 12768 32444 12774 32456
rect 13725 32453 13737 32456
rect 13771 32453 13783 32487
rect 13725 32447 13783 32453
rect 8849 32419 8907 32425
rect 8168 32388 8616 32416
rect 8168 32376 8174 32388
rect 7377 32351 7435 32357
rect 7377 32348 7389 32351
rect 5828 32320 7389 32348
rect 7377 32317 7389 32320
rect 7423 32348 7435 32351
rect 7466 32348 7472 32360
rect 7423 32320 7472 32348
rect 7423 32317 7435 32320
rect 7377 32311 7435 32317
rect 7466 32308 7472 32320
rect 7524 32308 7530 32360
rect 7561 32351 7619 32357
rect 7561 32317 7573 32351
rect 7607 32348 7619 32351
rect 8202 32348 8208 32360
rect 7607 32320 8208 32348
rect 7607 32317 7619 32320
rect 7561 32311 7619 32317
rect 8202 32308 8208 32320
rect 8260 32308 8266 32360
rect 8297 32351 8355 32357
rect 8297 32317 8309 32351
rect 8343 32348 8355 32351
rect 8386 32348 8392 32360
rect 8343 32320 8392 32348
rect 8343 32317 8355 32320
rect 8297 32311 8355 32317
rect 8386 32308 8392 32320
rect 8444 32308 8450 32360
rect 8588 32348 8616 32388
rect 8849 32385 8861 32419
rect 8895 32385 8907 32419
rect 11882 32416 11888 32428
rect 11843 32388 11888 32416
rect 8849 32379 8907 32385
rect 11882 32376 11888 32388
rect 11940 32376 11946 32428
rect 11977 32419 12035 32425
rect 11977 32385 11989 32419
rect 12023 32416 12035 32419
rect 12066 32416 12072 32428
rect 12023 32388 12072 32416
rect 12023 32385 12035 32388
rect 11977 32379 12035 32385
rect 12066 32376 12072 32388
rect 12124 32376 12130 32428
rect 12250 32416 12256 32428
rect 12211 32388 12256 32416
rect 12250 32376 12256 32388
rect 12308 32376 12314 32428
rect 8941 32351 8999 32357
rect 8941 32348 8953 32351
rect 8588 32320 8953 32348
rect 8941 32317 8953 32320
rect 8987 32317 8999 32351
rect 8941 32311 8999 32317
rect 12434 32308 12440 32360
rect 12492 32348 12498 32360
rect 12713 32351 12771 32357
rect 12713 32348 12725 32351
rect 12492 32320 12725 32348
rect 12492 32308 12498 32320
rect 12713 32317 12725 32320
rect 12759 32317 12771 32351
rect 12713 32311 12771 32317
rect 5813 32283 5871 32289
rect 5813 32249 5825 32283
rect 5859 32280 5871 32283
rect 7282 32280 7288 32292
rect 5859 32252 7288 32280
rect 5859 32249 5871 32252
rect 5813 32243 5871 32249
rect 7282 32240 7288 32252
rect 7340 32240 7346 32292
rect 11974 32240 11980 32292
rect 12032 32280 12038 32292
rect 12161 32283 12219 32289
rect 12161 32280 12173 32283
rect 12032 32252 12173 32280
rect 12032 32240 12038 32252
rect 12161 32249 12173 32252
rect 12207 32249 12219 32283
rect 12161 32243 12219 32249
rect 13081 32283 13139 32289
rect 13081 32249 13093 32283
rect 13127 32280 13139 32283
rect 13170 32280 13176 32292
rect 13127 32252 13176 32280
rect 13127 32249 13139 32252
rect 13081 32243 13139 32249
rect 13170 32240 13176 32252
rect 13228 32240 13234 32292
rect 4982 32212 4988 32224
rect 4943 32184 4988 32212
rect 4982 32172 4988 32184
rect 5040 32172 5046 32224
rect 6641 32215 6699 32221
rect 6641 32181 6653 32215
rect 6687 32212 6699 32215
rect 6914 32212 6920 32224
rect 6687 32184 6920 32212
rect 6687 32181 6699 32184
rect 6641 32175 6699 32181
rect 6914 32172 6920 32184
rect 6972 32172 6978 32224
rect 10870 32212 10876 32224
rect 10831 32184 10876 32212
rect 10870 32172 10876 32184
rect 10928 32212 10934 32224
rect 12342 32212 12348 32224
rect 10928 32184 12348 32212
rect 10928 32172 10934 32184
rect 12342 32172 12348 32184
rect 12400 32172 12406 32224
rect 13722 32172 13728 32224
rect 13780 32212 13786 32224
rect 13817 32215 13875 32221
rect 13817 32212 13829 32215
rect 13780 32184 13829 32212
rect 13780 32172 13786 32184
rect 13817 32181 13829 32184
rect 13863 32181 13875 32215
rect 13817 32175 13875 32181
rect 1104 32122 18860 32144
rect 1104 32070 3915 32122
rect 3967 32070 3979 32122
rect 4031 32070 4043 32122
rect 4095 32070 4107 32122
rect 4159 32070 4171 32122
rect 4223 32070 9846 32122
rect 9898 32070 9910 32122
rect 9962 32070 9974 32122
rect 10026 32070 10038 32122
rect 10090 32070 10102 32122
rect 10154 32070 15776 32122
rect 15828 32070 15840 32122
rect 15892 32070 15904 32122
rect 15956 32070 15968 32122
rect 16020 32070 16032 32122
rect 16084 32070 18860 32122
rect 1104 32048 18860 32070
rect 4246 32008 4252 32020
rect 4207 31980 4252 32008
rect 4246 31968 4252 31980
rect 4304 31968 4310 32020
rect 4522 31968 4528 32020
rect 4580 32008 4586 32020
rect 4801 32011 4859 32017
rect 4801 32008 4813 32011
rect 4580 31980 4813 32008
rect 4580 31968 4586 31980
rect 4801 31977 4813 31980
rect 4847 31977 4859 32011
rect 4801 31971 4859 31977
rect 5074 31968 5080 32020
rect 5132 32008 5138 32020
rect 5445 32011 5503 32017
rect 5445 32008 5457 32011
rect 5132 31980 5457 32008
rect 5132 31968 5138 31980
rect 5445 31977 5457 31980
rect 5491 31977 5503 32011
rect 5445 31971 5503 31977
rect 7466 31968 7472 32020
rect 7524 32008 7530 32020
rect 7745 32011 7803 32017
rect 7745 32008 7757 32011
rect 7524 31980 7757 32008
rect 7524 31968 7530 31980
rect 7745 31977 7757 31980
rect 7791 31977 7803 32011
rect 7745 31971 7803 31977
rect 9125 32011 9183 32017
rect 9125 31977 9137 32011
rect 9171 32008 9183 32011
rect 9582 32008 9588 32020
rect 9171 31980 9588 32008
rect 9171 31977 9183 31980
rect 9125 31971 9183 31977
rect 9582 31968 9588 31980
rect 9640 31968 9646 32020
rect 12618 31968 12624 32020
rect 12676 32008 12682 32020
rect 12713 32011 12771 32017
rect 12713 32008 12725 32011
rect 12676 31980 12725 32008
rect 12676 31968 12682 31980
rect 12713 31977 12725 31980
rect 12759 31977 12771 32011
rect 12713 31971 12771 31977
rect 7006 31940 7012 31952
rect 6104 31912 7012 31940
rect 3786 31832 3792 31884
rect 3844 31872 3850 31884
rect 3881 31875 3939 31881
rect 3881 31872 3893 31875
rect 3844 31844 3893 31872
rect 3844 31832 3850 31844
rect 3881 31841 3893 31844
rect 3927 31841 3939 31875
rect 5810 31872 5816 31884
rect 5771 31844 5816 31872
rect 3881 31835 3939 31841
rect 5810 31832 5816 31844
rect 5868 31832 5874 31884
rect 6104 31872 6132 31912
rect 7006 31900 7012 31912
rect 7064 31900 7070 31952
rect 7285 31943 7343 31949
rect 7285 31909 7297 31943
rect 7331 31909 7343 31943
rect 10965 31943 11023 31949
rect 10965 31940 10977 31943
rect 7285 31903 7343 31909
rect 9232 31912 10977 31940
rect 7300 31872 7328 31903
rect 9232 31881 9260 31912
rect 10965 31909 10977 31912
rect 11011 31909 11023 31943
rect 10965 31903 11023 31909
rect 5920 31844 6132 31872
rect 6196 31844 7328 31872
rect 9217 31875 9275 31881
rect 3970 31804 3976 31816
rect 3931 31776 3976 31804
rect 3970 31764 3976 31776
rect 4028 31764 4034 31816
rect 4798 31804 4804 31816
rect 4759 31776 4804 31804
rect 4798 31764 4804 31776
rect 4856 31764 4862 31816
rect 4982 31764 4988 31816
rect 5040 31804 5046 31816
rect 5626 31804 5632 31816
rect 5040 31776 5085 31804
rect 5587 31776 5632 31804
rect 5040 31764 5046 31776
rect 5626 31764 5632 31776
rect 5684 31764 5690 31816
rect 5718 31764 5724 31816
rect 5776 31804 5782 31816
rect 5920 31813 5948 31844
rect 5905 31807 5963 31813
rect 5905 31804 5917 31807
rect 5776 31776 5917 31804
rect 5776 31764 5782 31776
rect 5905 31773 5917 31776
rect 5951 31773 5963 31807
rect 5905 31767 5963 31773
rect 5997 31807 6055 31813
rect 5997 31773 6009 31807
rect 6043 31804 6055 31807
rect 6086 31804 6092 31816
rect 6043 31776 6092 31804
rect 6043 31773 6055 31776
rect 5997 31767 6055 31773
rect 6086 31764 6092 31776
rect 6144 31764 6150 31816
rect 6196 31813 6224 31844
rect 9217 31841 9229 31875
rect 9263 31841 9275 31875
rect 9217 31835 9275 31841
rect 9398 31832 9404 31884
rect 9456 31872 9462 31884
rect 10137 31875 10195 31881
rect 9456 31844 10088 31872
rect 9456 31832 9462 31844
rect 6181 31807 6239 31813
rect 6181 31773 6193 31807
rect 6227 31773 6239 31807
rect 6641 31807 6699 31813
rect 6641 31804 6653 31807
rect 6181 31767 6239 31773
rect 6288 31776 6653 31804
rect 5442 31696 5448 31748
rect 5500 31736 5506 31748
rect 6288 31736 6316 31776
rect 6641 31773 6653 31776
rect 6687 31773 6699 31807
rect 6641 31767 6699 31773
rect 6730 31764 6736 31816
rect 6788 31804 6794 31816
rect 7006 31804 7012 31816
rect 6788 31776 6833 31804
rect 6967 31776 7012 31804
rect 6788 31764 6794 31776
rect 7006 31764 7012 31776
rect 7064 31764 7070 31816
rect 7098 31764 7104 31816
rect 7156 31813 7162 31816
rect 7156 31804 7164 31813
rect 7926 31804 7932 31816
rect 7156 31776 7201 31804
rect 7887 31776 7932 31804
rect 7156 31767 7164 31776
rect 7156 31764 7162 31767
rect 7926 31764 7932 31776
rect 7984 31764 7990 31816
rect 10060 31813 10088 31844
rect 10137 31841 10149 31875
rect 10183 31872 10195 31875
rect 10318 31872 10324 31884
rect 10183 31844 10324 31872
rect 10183 31841 10195 31844
rect 10137 31835 10195 31841
rect 10318 31832 10324 31844
rect 10376 31832 10382 31884
rect 10410 31832 10416 31884
rect 10468 31872 10474 31884
rect 10468 31844 10732 31872
rect 10468 31832 10474 31844
rect 10704 31813 10732 31844
rect 10778 31832 10784 31884
rect 10836 31872 10842 31884
rect 11149 31875 11207 31881
rect 11149 31872 11161 31875
rect 10836 31844 11161 31872
rect 10836 31832 10842 31844
rect 11149 31841 11161 31844
rect 11195 31841 11207 31875
rect 11149 31835 11207 31841
rect 11701 31875 11759 31881
rect 11701 31841 11713 31875
rect 11747 31872 11759 31875
rect 12434 31872 12440 31884
rect 11747 31844 12440 31872
rect 11747 31841 11759 31844
rect 11701 31835 11759 31841
rect 12434 31832 12440 31844
rect 12492 31832 12498 31884
rect 8021 31807 8079 31813
rect 8021 31773 8033 31807
rect 8067 31804 8079 31807
rect 8941 31807 8999 31813
rect 8067 31776 8101 31804
rect 8067 31773 8079 31776
rect 8021 31767 8079 31773
rect 8941 31773 8953 31807
rect 8987 31773 8999 31807
rect 8941 31767 8999 31773
rect 9033 31807 9091 31813
rect 9033 31773 9045 31807
rect 9079 31804 9091 31807
rect 10045 31807 10103 31813
rect 9079 31776 9996 31804
rect 9079 31773 9091 31776
rect 9033 31767 9091 31773
rect 5500 31708 6316 31736
rect 5500 31696 5506 31708
rect 6914 31696 6920 31748
rect 6972 31736 6978 31748
rect 8036 31736 8064 31767
rect 6972 31708 7065 31736
rect 7852 31708 8064 31736
rect 6972 31696 6978 31708
rect 6932 31668 6960 31696
rect 7852 31680 7880 31708
rect 7834 31668 7840 31680
rect 6932 31640 7840 31668
rect 7834 31628 7840 31640
rect 7892 31628 7898 31680
rect 8956 31668 8984 31767
rect 9968 31736 9996 31776
rect 10045 31773 10057 31807
rect 10091 31804 10103 31807
rect 10689 31807 10747 31813
rect 10091 31776 10640 31804
rect 10091 31773 10103 31776
rect 10045 31767 10103 31773
rect 10410 31736 10416 31748
rect 9968 31708 10416 31736
rect 10410 31696 10416 31708
rect 10468 31696 10474 31748
rect 10612 31736 10640 31776
rect 10689 31773 10701 31807
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 11790 31764 11796 31816
rect 11848 31804 11854 31816
rect 11885 31807 11943 31813
rect 11885 31804 11897 31807
rect 11848 31776 11897 31804
rect 11848 31764 11854 31776
rect 11885 31773 11897 31776
rect 11931 31773 11943 31807
rect 11885 31767 11943 31773
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31804 12127 31807
rect 12529 31807 12587 31813
rect 12529 31804 12541 31807
rect 12115 31776 12541 31804
rect 12115 31773 12127 31776
rect 12069 31767 12127 31773
rect 12529 31773 12541 31776
rect 12575 31773 12587 31807
rect 12529 31767 12587 31773
rect 11146 31736 11152 31748
rect 10612 31708 11152 31736
rect 11146 31696 11152 31708
rect 11204 31696 11210 31748
rect 9677 31671 9735 31677
rect 9677 31668 9689 31671
rect 8956 31640 9689 31668
rect 9677 31637 9689 31640
rect 9723 31668 9735 31671
rect 9950 31668 9956 31680
rect 9723 31640 9956 31668
rect 9723 31637 9735 31640
rect 9677 31631 9735 31637
rect 9950 31628 9956 31640
rect 10008 31668 10014 31680
rect 10781 31671 10839 31677
rect 10781 31668 10793 31671
rect 10008 31640 10793 31668
rect 10008 31628 10014 31640
rect 10781 31637 10793 31640
rect 10827 31637 10839 31671
rect 10781 31631 10839 31637
rect 1104 31578 18860 31600
rect 1104 31526 6880 31578
rect 6932 31526 6944 31578
rect 6996 31526 7008 31578
rect 7060 31526 7072 31578
rect 7124 31526 7136 31578
rect 7188 31526 12811 31578
rect 12863 31526 12875 31578
rect 12927 31526 12939 31578
rect 12991 31526 13003 31578
rect 13055 31526 13067 31578
rect 13119 31526 18860 31578
rect 1104 31504 18860 31526
rect 2869 31467 2927 31473
rect 2869 31433 2881 31467
rect 2915 31464 2927 31467
rect 3050 31464 3056 31476
rect 2915 31436 3056 31464
rect 2915 31433 2927 31436
rect 2869 31427 2927 31433
rect 3050 31424 3056 31436
rect 3108 31464 3114 31476
rect 3970 31464 3976 31476
rect 3108 31436 3976 31464
rect 3108 31424 3114 31436
rect 3970 31424 3976 31436
rect 4028 31424 4034 31476
rect 5169 31467 5227 31473
rect 5169 31433 5181 31467
rect 5215 31464 5227 31467
rect 5626 31464 5632 31476
rect 5215 31436 5632 31464
rect 5215 31433 5227 31436
rect 5169 31427 5227 31433
rect 5626 31424 5632 31436
rect 5684 31464 5690 31476
rect 6730 31464 6736 31476
rect 5684 31436 6736 31464
rect 5684 31424 5690 31436
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 10134 31464 10140 31476
rect 9784 31436 10140 31464
rect 7282 31396 7288 31408
rect 2516 31368 4384 31396
rect 2516 31337 2544 31368
rect 4356 31337 4384 31368
rect 7024 31368 7288 31396
rect 2501 31331 2559 31337
rect 2501 31297 2513 31331
rect 2547 31297 2559 31331
rect 3513 31331 3571 31337
rect 3513 31328 3525 31331
rect 2501 31291 2559 31297
rect 2608 31300 3525 31328
rect 2608 31272 2636 31300
rect 3513 31297 3525 31300
rect 3559 31297 3571 31331
rect 3513 31291 3571 31297
rect 4341 31331 4399 31337
rect 4341 31297 4353 31331
rect 4387 31328 4399 31331
rect 4982 31328 4988 31340
rect 4387 31300 4988 31328
rect 4387 31297 4399 31300
rect 4341 31291 4399 31297
rect 4982 31288 4988 31300
rect 5040 31328 5046 31340
rect 7024 31337 7052 31368
rect 7282 31356 7288 31368
rect 7340 31356 7346 31408
rect 9122 31396 9128 31408
rect 8588 31368 9128 31396
rect 8588 31337 8616 31368
rect 9122 31356 9128 31368
rect 9180 31356 9186 31408
rect 5077 31331 5135 31337
rect 5077 31328 5089 31331
rect 5040 31300 5089 31328
rect 5040 31288 5046 31300
rect 5077 31297 5089 31300
rect 5123 31297 5135 31331
rect 5077 31291 5135 31297
rect 7009 31331 7067 31337
rect 7009 31297 7021 31331
rect 7055 31297 7067 31331
rect 7009 31291 7067 31297
rect 8573 31331 8631 31337
rect 8573 31297 8585 31331
rect 8619 31297 8631 31331
rect 8573 31291 8631 31297
rect 8665 31331 8723 31337
rect 8665 31297 8677 31331
rect 8711 31297 8723 31331
rect 8665 31291 8723 31297
rect 2590 31260 2596 31272
rect 2503 31232 2596 31260
rect 2590 31220 2596 31232
rect 2648 31220 2654 31272
rect 3329 31263 3387 31269
rect 3329 31229 3341 31263
rect 3375 31260 3387 31263
rect 3602 31260 3608 31272
rect 3375 31232 3608 31260
rect 3375 31229 3387 31232
rect 3329 31223 3387 31229
rect 3602 31220 3608 31232
rect 3660 31260 3666 31272
rect 4065 31263 4123 31269
rect 4065 31260 4077 31263
rect 3660 31232 4077 31260
rect 3660 31220 3666 31232
rect 4065 31229 4077 31232
rect 4111 31229 4123 31263
rect 4065 31223 4123 31229
rect 7285 31263 7343 31269
rect 7285 31229 7297 31263
rect 7331 31260 7343 31263
rect 7834 31260 7840 31272
rect 7331 31232 7840 31260
rect 7331 31229 7343 31232
rect 7285 31223 7343 31229
rect 7834 31220 7840 31232
rect 7892 31220 7898 31272
rect 8680 31192 8708 31291
rect 8754 31288 8760 31340
rect 8812 31328 8818 31340
rect 8941 31331 8999 31337
rect 8812 31300 8857 31328
rect 8812 31288 8818 31300
rect 8941 31297 8953 31331
rect 8987 31328 8999 31331
rect 9784 31328 9812 31436
rect 10134 31424 10140 31436
rect 10192 31424 10198 31476
rect 10321 31467 10379 31473
rect 10321 31433 10333 31467
rect 10367 31464 10379 31467
rect 10962 31464 10968 31476
rect 10367 31436 10968 31464
rect 10367 31433 10379 31436
rect 10321 31427 10379 31433
rect 10962 31424 10968 31436
rect 11020 31424 11026 31476
rect 11517 31399 11575 31405
rect 11517 31396 11529 31399
rect 9876 31368 11529 31396
rect 9876 31337 9904 31368
rect 11517 31365 11529 31368
rect 11563 31365 11575 31399
rect 11517 31359 11575 31365
rect 8987 31300 9812 31328
rect 9861 31331 9919 31337
rect 8987 31297 8999 31300
rect 8941 31291 8999 31297
rect 9861 31297 9873 31331
rect 9907 31297 9919 31331
rect 9861 31291 9919 31297
rect 9950 31288 9956 31340
rect 10008 31328 10014 31340
rect 10137 31331 10195 31337
rect 10008 31300 10053 31328
rect 10008 31288 10014 31300
rect 10137 31297 10149 31331
rect 10183 31297 10195 31331
rect 10137 31291 10195 31297
rect 8846 31220 8852 31272
rect 8904 31260 8910 31272
rect 9582 31260 9588 31272
rect 8904 31232 9588 31260
rect 8904 31220 8910 31232
rect 9582 31220 9588 31232
rect 9640 31260 9646 31272
rect 10152 31260 10180 31291
rect 10318 31288 10324 31340
rect 10376 31328 10382 31340
rect 10594 31328 10600 31340
rect 10376 31300 10600 31328
rect 10376 31288 10382 31300
rect 10594 31288 10600 31300
rect 10652 31288 10658 31340
rect 11146 31288 11152 31340
rect 11204 31328 11210 31340
rect 11793 31331 11851 31337
rect 11793 31328 11805 31331
rect 11204 31300 11805 31328
rect 11204 31288 11210 31300
rect 11793 31297 11805 31300
rect 11839 31297 11851 31331
rect 11793 31291 11851 31297
rect 14182 31288 14188 31340
rect 14240 31328 14246 31340
rect 14366 31328 14372 31340
rect 14240 31300 14372 31328
rect 14240 31288 14246 31300
rect 14366 31288 14372 31300
rect 14424 31288 14430 31340
rect 16850 31328 16856 31340
rect 16811 31300 16856 31328
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 9640 31232 10180 31260
rect 9640 31220 9646 31232
rect 10226 31220 10232 31272
rect 10284 31260 10290 31272
rect 11517 31263 11575 31269
rect 11517 31260 11529 31263
rect 10284 31232 11529 31260
rect 10284 31220 10290 31232
rect 11517 31229 11529 31232
rect 11563 31229 11575 31263
rect 11517 31223 11575 31229
rect 14274 31220 14280 31272
rect 14332 31260 14338 31272
rect 14553 31263 14611 31269
rect 14553 31260 14565 31263
rect 14332 31232 14565 31260
rect 14332 31220 14338 31232
rect 14553 31229 14565 31232
rect 14599 31229 14611 31263
rect 14553 31223 14611 31229
rect 9766 31192 9772 31204
rect 8680 31164 9772 31192
rect 9766 31152 9772 31164
rect 9824 31152 9830 31204
rect 10045 31195 10103 31201
rect 10045 31161 10057 31195
rect 10091 31192 10103 31195
rect 10594 31192 10600 31204
rect 10091 31164 10600 31192
rect 10091 31161 10103 31164
rect 10045 31155 10103 31161
rect 10594 31152 10600 31164
rect 10652 31152 10658 31204
rect 3510 31084 3516 31136
rect 3568 31124 3574 31136
rect 4157 31127 4215 31133
rect 4157 31124 4169 31127
rect 3568 31096 4169 31124
rect 3568 31084 3574 31096
rect 4157 31093 4169 31096
rect 4203 31093 4215 31127
rect 4157 31087 4215 31093
rect 4246 31084 4252 31136
rect 4304 31124 4310 31136
rect 6822 31124 6828 31136
rect 4304 31096 4349 31124
rect 6783 31096 6828 31124
rect 4304 31084 4310 31096
rect 6822 31084 6828 31096
rect 6880 31084 6886 31136
rect 7190 31124 7196 31136
rect 7151 31096 7196 31124
rect 7190 31084 7196 31096
rect 7248 31124 7254 31136
rect 7926 31124 7932 31136
rect 7248 31096 7932 31124
rect 7248 31084 7254 31096
rect 7926 31084 7932 31096
rect 7984 31084 7990 31136
rect 8294 31124 8300 31136
rect 8255 31096 8300 31124
rect 8294 31084 8300 31096
rect 8352 31084 8358 31136
rect 10962 31084 10968 31136
rect 11020 31124 11026 31136
rect 11701 31127 11759 31133
rect 11701 31124 11713 31127
rect 11020 31096 11713 31124
rect 11020 31084 11026 31096
rect 11701 31093 11713 31096
rect 11747 31093 11759 31127
rect 11701 31087 11759 31093
rect 13354 31084 13360 31136
rect 13412 31124 13418 31136
rect 14185 31127 14243 31133
rect 14185 31124 14197 31127
rect 13412 31096 14197 31124
rect 13412 31084 13418 31096
rect 14185 31093 14197 31096
rect 14231 31093 14243 31127
rect 16666 31124 16672 31136
rect 16627 31096 16672 31124
rect 14185 31087 14243 31093
rect 16666 31084 16672 31096
rect 16724 31084 16730 31136
rect 1104 31034 18860 31056
rect 1104 30982 3915 31034
rect 3967 30982 3979 31034
rect 4031 30982 4043 31034
rect 4095 30982 4107 31034
rect 4159 30982 4171 31034
rect 4223 30982 9846 31034
rect 9898 30982 9910 31034
rect 9962 30982 9974 31034
rect 10026 30982 10038 31034
rect 10090 30982 10102 31034
rect 10154 30982 15776 31034
rect 15828 30982 15840 31034
rect 15892 30982 15904 31034
rect 15956 30982 15968 31034
rect 16020 30982 16032 31034
rect 16084 30982 18860 31034
rect 1104 30960 18860 30982
rect 2682 30920 2688 30932
rect 2643 30892 2688 30920
rect 2682 30880 2688 30892
rect 2740 30880 2746 30932
rect 3786 30880 3792 30932
rect 3844 30920 3850 30932
rect 4065 30923 4123 30929
rect 4065 30920 4077 30923
rect 3844 30892 4077 30920
rect 3844 30880 3850 30892
rect 4065 30889 4077 30892
rect 4111 30889 4123 30923
rect 4065 30883 4123 30889
rect 8386 30880 8392 30932
rect 8444 30920 8450 30932
rect 9033 30923 9091 30929
rect 9033 30920 9045 30923
rect 8444 30892 9045 30920
rect 8444 30880 8450 30892
rect 9033 30889 9045 30892
rect 9079 30889 9091 30923
rect 9033 30883 9091 30889
rect 10410 30880 10416 30932
rect 10468 30920 10474 30932
rect 10689 30923 10747 30929
rect 10689 30920 10701 30923
rect 10468 30892 10701 30920
rect 10468 30880 10474 30892
rect 10689 30889 10701 30892
rect 10735 30889 10747 30923
rect 10689 30883 10747 30889
rect 3050 30852 3056 30864
rect 3011 30824 3056 30852
rect 3050 30812 3056 30824
rect 3108 30812 3114 30864
rect 10778 30784 10784 30796
rect 10739 30756 10784 30784
rect 10778 30744 10784 30756
rect 10836 30744 10842 30796
rect 2866 30716 2872 30728
rect 2827 30688 2872 30716
rect 2866 30676 2872 30688
rect 2924 30676 2930 30728
rect 2958 30676 2964 30728
rect 3016 30716 3022 30728
rect 3145 30719 3203 30725
rect 3016 30688 3061 30716
rect 3016 30676 3022 30688
rect 3145 30685 3157 30719
rect 3191 30716 3203 30719
rect 3510 30716 3516 30728
rect 3191 30688 3516 30716
rect 3191 30685 3203 30688
rect 3145 30679 3203 30685
rect 3510 30676 3516 30688
rect 3568 30676 3574 30728
rect 3602 30676 3608 30728
rect 3660 30716 3666 30728
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 3660 30688 3801 30716
rect 3660 30676 3666 30688
rect 3789 30685 3801 30688
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 6457 30719 6515 30725
rect 6457 30685 6469 30719
rect 6503 30716 6515 30719
rect 7282 30716 7288 30728
rect 6503 30688 7288 30716
rect 6503 30685 6515 30688
rect 6457 30679 6515 30685
rect 7282 30676 7288 30688
rect 7340 30676 7346 30728
rect 8941 30719 8999 30725
rect 8941 30685 8953 30719
rect 8987 30716 8999 30719
rect 9030 30716 9036 30728
rect 8987 30688 9036 30716
rect 8987 30685 8999 30688
rect 8941 30679 8999 30685
rect 9030 30676 9036 30688
rect 9088 30676 9094 30728
rect 9125 30719 9183 30725
rect 9125 30685 9137 30719
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 4065 30651 4123 30657
rect 4065 30648 4077 30651
rect 3804 30620 4077 30648
rect 3804 30592 3832 30620
rect 4065 30617 4077 30620
rect 4111 30617 4123 30651
rect 4065 30611 4123 30617
rect 6724 30651 6782 30657
rect 6724 30617 6736 30651
rect 6770 30648 6782 30651
rect 6822 30648 6828 30660
rect 6770 30620 6828 30648
rect 6770 30617 6782 30620
rect 6724 30611 6782 30617
rect 6822 30608 6828 30620
rect 6880 30608 6886 30660
rect 7190 30608 7196 30660
rect 7248 30648 7254 30660
rect 7374 30648 7380 30660
rect 7248 30620 7380 30648
rect 7248 30608 7254 30620
rect 7374 30608 7380 30620
rect 7432 30608 7438 30660
rect 7742 30608 7748 30660
rect 7800 30648 7806 30660
rect 9140 30648 9168 30679
rect 9582 30676 9588 30728
rect 9640 30716 9646 30728
rect 10505 30719 10563 30725
rect 10505 30716 10517 30719
rect 9640 30688 10517 30716
rect 9640 30676 9646 30688
rect 10505 30685 10517 30688
rect 10551 30685 10563 30719
rect 10505 30679 10563 30685
rect 10594 30676 10600 30728
rect 10652 30716 10658 30728
rect 13354 30716 13360 30728
rect 10652 30688 10697 30716
rect 13315 30688 13360 30716
rect 10652 30676 10658 30688
rect 13354 30676 13360 30688
rect 13412 30676 13418 30728
rect 15470 30716 15476 30728
rect 15431 30688 15476 30716
rect 15470 30676 15476 30688
rect 15528 30716 15534 30728
rect 17313 30719 17371 30725
rect 17313 30716 17325 30719
rect 15528 30688 17325 30716
rect 15528 30676 15534 30688
rect 17313 30685 17325 30688
rect 17359 30685 17371 30719
rect 17313 30679 17371 30685
rect 9674 30648 9680 30660
rect 7800 30620 9076 30648
rect 9140 30620 9680 30648
rect 7800 30608 7806 30620
rect 3786 30540 3792 30592
rect 3844 30540 3850 30592
rect 3881 30583 3939 30589
rect 3881 30549 3893 30583
rect 3927 30580 3939 30583
rect 4246 30580 4252 30592
rect 3927 30552 4252 30580
rect 3927 30549 3939 30552
rect 3881 30543 3939 30549
rect 4246 30540 4252 30552
rect 4304 30540 4310 30592
rect 7834 30580 7840 30592
rect 7795 30552 7840 30580
rect 7834 30540 7840 30552
rect 7892 30540 7898 30592
rect 9048 30580 9076 30620
rect 9674 30608 9680 30620
rect 9732 30608 9738 30660
rect 9861 30651 9919 30657
rect 9861 30617 9873 30651
rect 9907 30648 9919 30651
rect 10962 30648 10968 30660
rect 9907 30620 10968 30648
rect 9907 30617 9919 30620
rect 9861 30611 9919 30617
rect 9876 30580 9904 30611
rect 10962 30608 10968 30620
rect 11020 30608 11026 30660
rect 15228 30651 15286 30657
rect 15228 30617 15240 30651
rect 15274 30648 15286 30651
rect 15746 30648 15752 30660
rect 15274 30620 15752 30648
rect 15274 30617 15286 30620
rect 15228 30611 15286 30617
rect 15746 30608 15752 30620
rect 15804 30608 15810 30660
rect 17068 30651 17126 30657
rect 17068 30617 17080 30651
rect 17114 30648 17126 30651
rect 17494 30648 17500 30660
rect 17114 30620 17500 30648
rect 17114 30617 17126 30620
rect 17068 30611 17126 30617
rect 17494 30608 17500 30620
rect 17552 30608 17558 30660
rect 9950 30580 9956 30592
rect 9048 30552 9956 30580
rect 9950 30540 9956 30552
rect 10008 30540 10014 30592
rect 10045 30583 10103 30589
rect 10045 30549 10057 30583
rect 10091 30580 10103 30583
rect 10410 30580 10416 30592
rect 10091 30552 10416 30580
rect 10091 30549 10103 30552
rect 10045 30543 10103 30549
rect 10410 30540 10416 30552
rect 10468 30540 10474 30592
rect 13541 30583 13599 30589
rect 13541 30549 13553 30583
rect 13587 30580 13599 30583
rect 13998 30580 14004 30592
rect 13587 30552 14004 30580
rect 13587 30549 13599 30552
rect 13541 30543 13599 30549
rect 13998 30540 14004 30552
rect 14056 30540 14062 30592
rect 14093 30583 14151 30589
rect 14093 30549 14105 30583
rect 14139 30580 14151 30583
rect 14274 30580 14280 30592
rect 14139 30552 14280 30580
rect 14139 30549 14151 30552
rect 14093 30543 14151 30549
rect 14274 30540 14280 30552
rect 14332 30540 14338 30592
rect 15933 30583 15991 30589
rect 15933 30549 15945 30583
rect 15979 30580 15991 30583
rect 16574 30580 16580 30592
rect 15979 30552 16580 30580
rect 15979 30549 15991 30552
rect 15933 30543 15991 30549
rect 16574 30540 16580 30552
rect 16632 30540 16638 30592
rect 1104 30490 18860 30512
rect 1104 30438 6880 30490
rect 6932 30438 6944 30490
rect 6996 30438 7008 30490
rect 7060 30438 7072 30490
rect 7124 30438 7136 30490
rect 7188 30438 12811 30490
rect 12863 30438 12875 30490
rect 12927 30438 12939 30490
rect 12991 30438 13003 30490
rect 13055 30438 13067 30490
rect 13119 30438 18860 30490
rect 1104 30416 18860 30438
rect 9030 30336 9036 30388
rect 9088 30376 9094 30388
rect 9125 30379 9183 30385
rect 9125 30376 9137 30379
rect 9088 30348 9137 30376
rect 9088 30336 9094 30348
rect 9125 30345 9137 30348
rect 9171 30345 9183 30379
rect 15746 30376 15752 30388
rect 15707 30348 15752 30376
rect 9125 30339 9183 30345
rect 15746 30336 15752 30348
rect 15804 30336 15810 30388
rect 16669 30379 16727 30385
rect 16669 30345 16681 30379
rect 16715 30376 16727 30379
rect 16850 30376 16856 30388
rect 16715 30348 16856 30376
rect 16715 30345 16727 30348
rect 16669 30339 16727 30345
rect 16850 30336 16856 30348
rect 16908 30336 16914 30388
rect 17494 30376 17500 30388
rect 17455 30348 17500 30376
rect 17494 30336 17500 30348
rect 17552 30336 17558 30388
rect 8012 30311 8070 30317
rect 8012 30277 8024 30311
rect 8058 30308 8070 30311
rect 8294 30308 8300 30320
rect 8058 30280 8300 30308
rect 8058 30277 8070 30280
rect 8012 30271 8070 30277
rect 8294 30268 8300 30280
rect 8352 30268 8358 30320
rect 9950 30268 9956 30320
rect 10008 30308 10014 30320
rect 15470 30308 15476 30320
rect 10008 30280 10088 30308
rect 10008 30268 10014 30280
rect 7282 30200 7288 30252
rect 7340 30240 7346 30252
rect 7745 30243 7803 30249
rect 7745 30240 7757 30243
rect 7340 30212 7757 30240
rect 7340 30200 7346 30212
rect 7745 30209 7757 30212
rect 7791 30209 7803 30243
rect 7745 30203 7803 30209
rect 9674 30200 9680 30252
rect 9732 30240 9738 30252
rect 10060 30249 10088 30280
rect 13924 30280 15476 30308
rect 9861 30243 9919 30249
rect 9861 30240 9873 30243
rect 9732 30212 9873 30240
rect 9732 30200 9738 30212
rect 9861 30209 9873 30212
rect 9907 30209 9919 30243
rect 9861 30203 9919 30209
rect 10045 30243 10103 30249
rect 10045 30209 10057 30243
rect 10091 30240 10103 30243
rect 10226 30240 10232 30252
rect 10091 30212 10232 30240
rect 10091 30209 10103 30212
rect 10045 30203 10103 30209
rect 10226 30200 10232 30212
rect 10284 30200 10290 30252
rect 10410 30200 10416 30252
rect 10468 30240 10474 30252
rect 10505 30243 10563 30249
rect 10505 30240 10517 30243
rect 10468 30212 10517 30240
rect 10468 30200 10474 30212
rect 10505 30209 10517 30212
rect 10551 30209 10563 30243
rect 10505 30203 10563 30209
rect 10689 30243 10747 30249
rect 10689 30209 10701 30243
rect 10735 30240 10747 30243
rect 10778 30240 10784 30252
rect 10735 30212 10784 30240
rect 10735 30209 10747 30212
rect 10689 30203 10747 30209
rect 9953 30175 10011 30181
rect 9953 30141 9965 30175
rect 9999 30172 10011 30175
rect 10704 30172 10732 30203
rect 10778 30200 10784 30212
rect 10836 30200 10842 30252
rect 13722 30240 13728 30252
rect 12406 30212 13728 30240
rect 9999 30144 10732 30172
rect 9999 30141 10011 30144
rect 9953 30135 10011 30141
rect 11330 30132 11336 30184
rect 11388 30172 11394 30184
rect 12406 30172 12434 30212
rect 13722 30200 13728 30212
rect 13780 30240 13786 30252
rect 13924 30249 13952 30280
rect 15470 30268 15476 30280
rect 15528 30268 15534 30320
rect 13909 30243 13967 30249
rect 13909 30240 13921 30243
rect 13780 30212 13921 30240
rect 13780 30200 13786 30212
rect 13909 30209 13921 30212
rect 13955 30209 13967 30243
rect 13909 30203 13967 30209
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 14165 30243 14223 30249
rect 14165 30240 14177 30243
rect 14056 30212 14177 30240
rect 14056 30200 14062 30212
rect 14165 30209 14177 30212
rect 14211 30209 14223 30243
rect 14165 30203 14223 30209
rect 14458 30200 14464 30252
rect 14516 30240 14522 30252
rect 15933 30243 15991 30249
rect 15933 30240 15945 30243
rect 14516 30212 15945 30240
rect 14516 30200 14522 30212
rect 15933 30209 15945 30212
rect 15979 30209 15991 30243
rect 15933 30203 15991 30209
rect 16758 30200 16764 30252
rect 16816 30240 16822 30252
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 16816 30212 16865 30240
rect 16816 30200 16822 30212
rect 16853 30209 16865 30212
rect 16899 30240 16911 30243
rect 16942 30240 16948 30252
rect 16899 30212 16948 30240
rect 16899 30209 16911 30212
rect 16853 30203 16911 30209
rect 16942 30200 16948 30212
rect 17000 30200 17006 30252
rect 17678 30240 17684 30252
rect 17639 30212 17684 30240
rect 17678 30200 17684 30212
rect 17736 30200 17742 30252
rect 11388 30144 12434 30172
rect 11388 30132 11394 30144
rect 16574 30132 16580 30184
rect 16632 30172 16638 30184
rect 17037 30175 17095 30181
rect 17037 30172 17049 30175
rect 16632 30144 17049 30172
rect 16632 30132 16638 30144
rect 17037 30141 17049 30144
rect 17083 30141 17095 30175
rect 17037 30135 17095 30141
rect 9674 29996 9680 30048
rect 9732 30036 9738 30048
rect 10594 30036 10600 30048
rect 9732 30008 10600 30036
rect 9732 29996 9738 30008
rect 10594 29996 10600 30008
rect 10652 29996 10658 30048
rect 15102 29996 15108 30048
rect 15160 30036 15166 30048
rect 15289 30039 15347 30045
rect 15289 30036 15301 30039
rect 15160 30008 15301 30036
rect 15160 29996 15166 30008
rect 15289 30005 15301 30008
rect 15335 30005 15347 30039
rect 15289 29999 15347 30005
rect 1104 29946 18860 29968
rect 1104 29894 3915 29946
rect 3967 29894 3979 29946
rect 4031 29894 4043 29946
rect 4095 29894 4107 29946
rect 4159 29894 4171 29946
rect 4223 29894 9846 29946
rect 9898 29894 9910 29946
rect 9962 29894 9974 29946
rect 10026 29894 10038 29946
rect 10090 29894 10102 29946
rect 10154 29894 15776 29946
rect 15828 29894 15840 29946
rect 15892 29894 15904 29946
rect 15956 29894 15968 29946
rect 16020 29894 16032 29946
rect 16084 29894 18860 29946
rect 1104 29872 18860 29894
rect 5442 29832 5448 29844
rect 5403 29804 5448 29832
rect 5442 29792 5448 29804
rect 5500 29792 5506 29844
rect 12526 29792 12532 29844
rect 12584 29832 12590 29844
rect 12713 29835 12771 29841
rect 12713 29832 12725 29835
rect 12584 29804 12725 29832
rect 12584 29792 12590 29804
rect 12713 29801 12725 29804
rect 12759 29801 12771 29835
rect 13722 29832 13728 29844
rect 12713 29795 12771 29801
rect 13188 29804 13728 29832
rect 3237 29767 3295 29773
rect 3237 29733 3249 29767
rect 3283 29764 3295 29767
rect 3786 29764 3792 29776
rect 3283 29736 3792 29764
rect 3283 29733 3295 29736
rect 3237 29727 3295 29733
rect 3786 29724 3792 29736
rect 3844 29724 3850 29776
rect 2958 29656 2964 29708
rect 3016 29696 3022 29708
rect 5813 29699 5871 29705
rect 3016 29668 3280 29696
rect 3016 29656 3022 29668
rect 2866 29588 2872 29640
rect 2924 29628 2930 29640
rect 3252 29637 3280 29668
rect 5813 29665 5825 29699
rect 5859 29696 5871 29699
rect 7834 29696 7840 29708
rect 5859 29668 7840 29696
rect 5859 29665 5871 29668
rect 5813 29659 5871 29665
rect 7834 29656 7840 29668
rect 7892 29656 7898 29708
rect 9674 29696 9680 29708
rect 9635 29668 9680 29696
rect 9674 29656 9680 29668
rect 9732 29656 9738 29708
rect 13188 29705 13216 29804
rect 13722 29792 13728 29804
rect 13780 29832 13786 29844
rect 14277 29835 14335 29841
rect 14277 29832 14289 29835
rect 13780 29804 14289 29832
rect 13780 29792 13786 29804
rect 14277 29801 14289 29804
rect 14323 29801 14335 29835
rect 14277 29795 14335 29801
rect 13541 29767 13599 29773
rect 13541 29733 13553 29767
rect 13587 29764 13599 29767
rect 14458 29764 14464 29776
rect 13587 29736 14464 29764
rect 13587 29733 13599 29736
rect 13541 29727 13599 29733
rect 14458 29724 14464 29736
rect 14516 29724 14522 29776
rect 13173 29699 13231 29705
rect 13173 29665 13185 29699
rect 13219 29665 13231 29699
rect 14182 29696 14188 29708
rect 13173 29659 13231 29665
rect 13372 29668 14188 29696
rect 13372 29640 13400 29668
rect 14182 29656 14188 29668
rect 14240 29696 14246 29708
rect 14240 29668 15240 29696
rect 14240 29656 14246 29668
rect 3053 29631 3111 29637
rect 3053 29628 3065 29631
rect 2924 29600 3065 29628
rect 2924 29588 2930 29600
rect 3053 29597 3065 29600
rect 3099 29597 3111 29631
rect 3053 29591 3111 29597
rect 3237 29631 3295 29637
rect 3237 29597 3249 29631
rect 3283 29597 3295 29631
rect 5626 29628 5632 29640
rect 5587 29600 5632 29628
rect 3237 29591 3295 29597
rect 5626 29588 5632 29600
rect 5684 29588 5690 29640
rect 5902 29628 5908 29640
rect 5863 29600 5908 29628
rect 5902 29588 5908 29600
rect 5960 29588 5966 29640
rect 5997 29631 6055 29637
rect 5997 29597 6009 29631
rect 6043 29628 6055 29631
rect 6086 29628 6092 29640
rect 6043 29600 6092 29628
rect 6043 29597 6055 29600
rect 5997 29591 6055 29597
rect 6086 29588 6092 29600
rect 6144 29588 6150 29640
rect 6181 29631 6239 29637
rect 6181 29597 6193 29631
rect 6227 29628 6239 29631
rect 6270 29628 6276 29640
rect 6227 29600 6276 29628
rect 6227 29597 6239 29600
rect 6181 29591 6239 29597
rect 6270 29588 6276 29600
rect 6328 29588 6334 29640
rect 9582 29628 9588 29640
rect 9543 29600 9588 29628
rect 9582 29588 9588 29600
rect 9640 29588 9646 29640
rect 10226 29588 10232 29640
rect 10284 29588 10290 29640
rect 11330 29628 11336 29640
rect 11291 29600 11336 29628
rect 11330 29588 11336 29600
rect 11388 29588 11394 29640
rect 13354 29628 13360 29640
rect 13315 29600 13360 29628
rect 13354 29588 13360 29600
rect 13412 29588 13418 29640
rect 14274 29628 14280 29640
rect 14235 29600 14280 29628
rect 14274 29588 14280 29600
rect 14332 29588 14338 29640
rect 14366 29588 14372 29640
rect 14424 29628 14430 29640
rect 15013 29631 15071 29637
rect 14424 29600 14469 29628
rect 14424 29588 14430 29600
rect 15013 29597 15025 29631
rect 15059 29628 15071 29631
rect 15102 29628 15108 29640
rect 15059 29600 15108 29628
rect 15059 29597 15071 29600
rect 15013 29591 15071 29597
rect 9674 29520 9680 29572
rect 9732 29560 9738 29572
rect 10244 29560 10272 29588
rect 9732 29532 10272 29560
rect 11600 29563 11658 29569
rect 9732 29520 9738 29532
rect 11600 29529 11612 29563
rect 11646 29560 11658 29563
rect 12066 29560 12072 29572
rect 11646 29532 12072 29560
rect 11646 29529 11658 29532
rect 11600 29523 11658 29529
rect 12066 29520 12072 29532
rect 12124 29520 12130 29572
rect 14550 29560 14556 29572
rect 14511 29532 14556 29560
rect 14550 29520 14556 29532
rect 14608 29560 14614 29572
rect 15028 29560 15056 29591
rect 15102 29588 15108 29600
rect 15160 29588 15166 29640
rect 15212 29637 15240 29668
rect 15470 29656 15476 29708
rect 15528 29696 15534 29708
rect 16209 29699 16267 29705
rect 16209 29696 16221 29699
rect 15528 29668 16221 29696
rect 15528 29656 15534 29668
rect 16209 29665 16221 29668
rect 16255 29665 16267 29699
rect 16209 29659 16267 29665
rect 15197 29631 15255 29637
rect 15197 29597 15209 29631
rect 15243 29597 15255 29631
rect 15197 29591 15255 29597
rect 14608 29532 15056 29560
rect 16476 29563 16534 29569
rect 14608 29520 14614 29532
rect 16476 29529 16488 29563
rect 16522 29560 16534 29563
rect 16666 29560 16672 29572
rect 16522 29532 16672 29560
rect 16522 29529 16534 29532
rect 16476 29523 16534 29529
rect 16666 29520 16672 29532
rect 16724 29520 16730 29572
rect 9953 29495 10011 29501
rect 9953 29461 9965 29495
rect 9999 29492 10011 29495
rect 10226 29492 10232 29504
rect 9999 29464 10232 29492
rect 9999 29461 10011 29464
rect 9953 29455 10011 29461
rect 10226 29452 10232 29464
rect 10284 29452 10290 29504
rect 13630 29452 13636 29504
rect 13688 29492 13694 29504
rect 14093 29495 14151 29501
rect 14093 29492 14105 29495
rect 13688 29464 14105 29492
rect 13688 29452 13694 29464
rect 14093 29461 14105 29464
rect 14139 29461 14151 29495
rect 14093 29455 14151 29461
rect 15381 29495 15439 29501
rect 15381 29461 15393 29495
rect 15427 29492 15439 29495
rect 15838 29492 15844 29504
rect 15427 29464 15844 29492
rect 15427 29461 15439 29464
rect 15381 29455 15439 29461
rect 15838 29452 15844 29464
rect 15896 29452 15902 29504
rect 17586 29492 17592 29504
rect 17547 29464 17592 29492
rect 17586 29452 17592 29464
rect 17644 29452 17650 29504
rect 1104 29402 18860 29424
rect 1104 29350 6880 29402
rect 6932 29350 6944 29402
rect 6996 29350 7008 29402
rect 7060 29350 7072 29402
rect 7124 29350 7136 29402
rect 7188 29350 12811 29402
rect 12863 29350 12875 29402
rect 12927 29350 12939 29402
rect 12991 29350 13003 29402
rect 13055 29350 13067 29402
rect 13119 29350 18860 29402
rect 1104 29328 18860 29350
rect 2869 29291 2927 29297
rect 2869 29257 2881 29291
rect 2915 29288 2927 29291
rect 2958 29288 2964 29300
rect 2915 29260 2964 29288
rect 2915 29257 2927 29260
rect 2869 29251 2927 29257
rect 2958 29248 2964 29260
rect 3016 29248 3022 29300
rect 5169 29291 5227 29297
rect 5169 29257 5181 29291
rect 5215 29288 5227 29291
rect 5902 29288 5908 29300
rect 5215 29260 5908 29288
rect 5215 29257 5227 29260
rect 5169 29251 5227 29257
rect 5902 29248 5908 29260
rect 5960 29248 5966 29300
rect 13817 29291 13875 29297
rect 13817 29257 13829 29291
rect 13863 29288 13875 29291
rect 14366 29288 14372 29300
rect 13863 29260 14372 29288
rect 13863 29257 13875 29260
rect 13817 29251 13875 29257
rect 14366 29248 14372 29260
rect 14424 29248 14430 29300
rect 15657 29291 15715 29297
rect 15657 29257 15669 29291
rect 15703 29257 15715 29291
rect 15657 29251 15715 29257
rect 17037 29291 17095 29297
rect 17037 29257 17049 29291
rect 17083 29288 17095 29291
rect 17678 29288 17684 29300
rect 17083 29260 17684 29288
rect 17083 29257 17095 29260
rect 17037 29251 17095 29257
rect 2501 29155 2559 29161
rect 2501 29121 2513 29155
rect 2547 29152 2559 29155
rect 2976 29152 3004 29248
rect 14952 29223 15010 29229
rect 14952 29189 14964 29223
rect 14998 29220 15010 29223
rect 15672 29220 15700 29251
rect 17678 29248 17684 29260
rect 17736 29248 17742 29300
rect 14998 29192 15700 29220
rect 14998 29189 15010 29192
rect 14952 29183 15010 29189
rect 3513 29155 3571 29161
rect 3513 29152 3525 29155
rect 2547 29124 2820 29152
rect 2976 29124 3525 29152
rect 2547 29121 2559 29124
rect 2501 29115 2559 29121
rect 2590 29084 2596 29096
rect 2551 29056 2596 29084
rect 2590 29044 2596 29056
rect 2648 29044 2654 29096
rect 2792 29016 2820 29124
rect 3513 29121 3525 29124
rect 3559 29121 3571 29155
rect 3513 29115 3571 29121
rect 3786 29112 3792 29164
rect 3844 29152 3850 29164
rect 4157 29155 4215 29161
rect 4157 29152 4169 29155
rect 3844 29124 4169 29152
rect 3844 29112 3850 29124
rect 4157 29121 4169 29124
rect 4203 29121 4215 29155
rect 4157 29115 4215 29121
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29121 5135 29155
rect 5077 29115 5135 29121
rect 15197 29155 15255 29161
rect 15197 29121 15209 29155
rect 15243 29152 15255 29155
rect 15470 29152 15476 29164
rect 15243 29124 15476 29152
rect 15243 29121 15255 29124
rect 15197 29115 15255 29121
rect 2866 29044 2872 29096
rect 2924 29084 2930 29096
rect 3326 29084 3332 29096
rect 2924 29056 3332 29084
rect 2924 29044 2930 29056
rect 3326 29044 3332 29056
rect 3384 29044 3390 29096
rect 3697 29087 3755 29093
rect 3697 29053 3709 29087
rect 3743 29084 3755 29087
rect 4249 29087 4307 29093
rect 4249 29084 4261 29087
rect 3743 29056 4261 29084
rect 3743 29053 3755 29056
rect 3697 29047 3755 29053
rect 4249 29053 4261 29056
rect 4295 29053 4307 29087
rect 4249 29047 4307 29053
rect 4433 29087 4491 29093
rect 4433 29053 4445 29087
rect 4479 29084 4491 29087
rect 4798 29084 4804 29096
rect 4479 29056 4804 29084
rect 4479 29053 4491 29056
rect 4433 29047 4491 29053
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 4154 29016 4160 29028
rect 2792 28988 4160 29016
rect 4154 28976 4160 28988
rect 4212 29016 4218 29028
rect 5092 29016 5120 29115
rect 15470 29112 15476 29124
rect 15528 29112 15534 29164
rect 15838 29152 15844 29164
rect 15799 29124 15844 29152
rect 15838 29112 15844 29124
rect 15896 29112 15902 29164
rect 16758 29152 16764 29164
rect 16719 29124 16764 29152
rect 16758 29112 16764 29124
rect 16816 29112 16822 29164
rect 16853 29155 16911 29161
rect 16853 29121 16865 29155
rect 16899 29152 16911 29155
rect 16942 29152 16948 29164
rect 16899 29124 16948 29152
rect 16899 29121 16911 29124
rect 16853 29115 16911 29121
rect 16942 29112 16948 29124
rect 17000 29112 17006 29164
rect 5258 29016 5264 29028
rect 4212 28988 5264 29016
rect 4212 28976 4218 28988
rect 5258 28976 5264 28988
rect 5316 28976 5322 29028
rect 4246 28908 4252 28960
rect 4304 28948 4310 28960
rect 4341 28951 4399 28957
rect 4341 28948 4353 28951
rect 4304 28920 4353 28948
rect 4304 28908 4310 28920
rect 4341 28917 4353 28920
rect 4387 28917 4399 28951
rect 4341 28911 4399 28917
rect 1104 28858 18860 28880
rect 1104 28806 3915 28858
rect 3967 28806 3979 28858
rect 4031 28806 4043 28858
rect 4095 28806 4107 28858
rect 4159 28806 4171 28858
rect 4223 28806 9846 28858
rect 9898 28806 9910 28858
rect 9962 28806 9974 28858
rect 10026 28806 10038 28858
rect 10090 28806 10102 28858
rect 10154 28806 15776 28858
rect 15828 28806 15840 28858
rect 15892 28806 15904 28858
rect 15956 28806 15968 28858
rect 16020 28806 16032 28858
rect 16084 28806 18860 28858
rect 1104 28784 18860 28806
rect 6270 28744 6276 28756
rect 6231 28716 6276 28744
rect 6270 28704 6276 28716
rect 6328 28704 6334 28756
rect 12066 28744 12072 28756
rect 12027 28716 12072 28744
rect 12066 28704 12072 28716
rect 12124 28704 12130 28756
rect 16758 28704 16764 28756
rect 16816 28744 16822 28756
rect 17129 28747 17187 28753
rect 17129 28744 17141 28747
rect 16816 28716 17141 28744
rect 16816 28704 16822 28716
rect 17129 28713 17141 28716
rect 17175 28713 17187 28747
rect 17129 28707 17187 28713
rect 14274 28636 14280 28688
rect 14332 28676 14338 28688
rect 14645 28679 14703 28685
rect 14645 28676 14657 28679
rect 14332 28648 14657 28676
rect 14332 28636 14338 28648
rect 14645 28645 14657 28648
rect 14691 28645 14703 28679
rect 14645 28639 14703 28645
rect 5902 28568 5908 28620
rect 5960 28608 5966 28620
rect 12437 28611 12495 28617
rect 5960 28580 6040 28608
rect 5960 28568 5966 28580
rect 3602 28500 3608 28552
rect 3660 28540 3666 28552
rect 3881 28543 3939 28549
rect 3881 28540 3893 28543
rect 3660 28512 3893 28540
rect 3660 28500 3666 28512
rect 3881 28509 3893 28512
rect 3927 28509 3939 28543
rect 3881 28503 3939 28509
rect 5534 28500 5540 28552
rect 5592 28540 5598 28552
rect 6012 28549 6040 28580
rect 12437 28577 12449 28611
rect 12483 28608 12495 28611
rect 12618 28608 12624 28620
rect 12483 28580 12624 28608
rect 12483 28577 12495 28580
rect 12437 28571 12495 28577
rect 12618 28568 12624 28580
rect 12676 28608 12682 28620
rect 13081 28611 13139 28617
rect 13081 28608 13093 28611
rect 12676 28580 13093 28608
rect 12676 28568 12682 28580
rect 13081 28577 13093 28580
rect 13127 28577 13139 28611
rect 13081 28571 13139 28577
rect 13722 28568 13728 28620
rect 13780 28608 13786 28620
rect 13780 28580 14504 28608
rect 13780 28568 13786 28580
rect 5721 28543 5779 28549
rect 5721 28540 5733 28543
rect 5592 28512 5733 28540
rect 5592 28500 5598 28512
rect 5721 28509 5733 28512
rect 5767 28509 5779 28543
rect 5721 28503 5779 28509
rect 5997 28543 6055 28549
rect 5997 28509 6009 28543
rect 6043 28509 6055 28543
rect 5997 28503 6055 28509
rect 6086 28500 6092 28552
rect 6144 28540 6150 28552
rect 7285 28543 7343 28549
rect 6144 28512 6189 28540
rect 6144 28500 6150 28512
rect 7285 28509 7297 28543
rect 7331 28540 7343 28543
rect 7374 28540 7380 28552
rect 7331 28512 7380 28540
rect 7331 28509 7343 28512
rect 7285 28503 7343 28509
rect 7374 28500 7380 28512
rect 7432 28500 7438 28552
rect 7469 28543 7527 28549
rect 7469 28509 7481 28543
rect 7515 28540 7527 28543
rect 7834 28540 7840 28552
rect 7515 28512 7840 28540
rect 7515 28509 7527 28512
rect 7469 28503 7527 28509
rect 7834 28500 7840 28512
rect 7892 28500 7898 28552
rect 10137 28543 10195 28549
rect 10137 28509 10149 28543
rect 10183 28540 10195 28543
rect 10226 28540 10232 28552
rect 10183 28512 10232 28540
rect 10183 28509 10195 28512
rect 10137 28503 10195 28509
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 10321 28543 10379 28549
rect 10321 28509 10333 28543
rect 10367 28540 10379 28543
rect 10870 28540 10876 28552
rect 10367 28512 10876 28540
rect 10367 28509 10379 28512
rect 10321 28503 10379 28509
rect 10870 28500 10876 28512
rect 10928 28500 10934 28552
rect 12253 28543 12311 28549
rect 12253 28509 12265 28543
rect 12299 28509 12311 28543
rect 12253 28503 12311 28509
rect 3786 28432 3792 28484
rect 3844 28472 3850 28484
rect 4126 28475 4184 28481
rect 4126 28472 4138 28475
rect 3844 28444 4138 28472
rect 3844 28432 3850 28444
rect 4126 28441 4138 28444
rect 4172 28441 4184 28475
rect 5902 28472 5908 28484
rect 5863 28444 5908 28472
rect 4126 28435 4184 28441
rect 5902 28432 5908 28444
rect 5960 28432 5966 28484
rect 12268 28472 12296 28503
rect 12342 28500 12348 28552
rect 12400 28540 12406 28552
rect 12529 28543 12587 28549
rect 12400 28512 12445 28540
rect 12400 28500 12406 28512
rect 12529 28509 12541 28543
rect 12575 28540 12587 28543
rect 12710 28540 12716 28552
rect 12575 28512 12716 28540
rect 12575 28509 12587 28512
rect 12529 28503 12587 28509
rect 12710 28500 12716 28512
rect 12768 28500 12774 28552
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28540 13323 28543
rect 13354 28540 13360 28552
rect 13311 28512 13360 28540
rect 13311 28509 13323 28512
rect 13265 28503 13323 28509
rect 13354 28500 13360 28512
rect 13412 28500 13418 28552
rect 14366 28540 14372 28552
rect 14327 28512 14372 28540
rect 14366 28500 14372 28512
rect 14424 28500 14430 28552
rect 14476 28549 14504 28580
rect 15470 28568 15476 28620
rect 15528 28608 15534 28620
rect 15749 28611 15807 28617
rect 15749 28608 15761 28611
rect 15528 28580 15761 28608
rect 15528 28568 15534 28580
rect 15749 28577 15761 28580
rect 15795 28577 15807 28611
rect 15749 28571 15807 28577
rect 14461 28543 14519 28549
rect 14461 28509 14473 28543
rect 14507 28509 14519 28543
rect 14461 28503 14519 28509
rect 13538 28472 13544 28484
rect 12268 28444 13544 28472
rect 13538 28432 13544 28444
rect 13596 28432 13602 28484
rect 13814 28432 13820 28484
rect 13872 28472 13878 28484
rect 14093 28475 14151 28481
rect 14093 28472 14105 28475
rect 13872 28444 14105 28472
rect 13872 28432 13878 28444
rect 14093 28441 14105 28444
rect 14139 28441 14151 28475
rect 14093 28435 14151 28441
rect 14277 28475 14335 28481
rect 14277 28441 14289 28475
rect 14323 28472 14335 28475
rect 14550 28472 14556 28484
rect 14323 28444 14556 28472
rect 14323 28441 14335 28444
rect 14277 28435 14335 28441
rect 14550 28432 14556 28444
rect 14608 28432 14614 28484
rect 16016 28475 16074 28481
rect 16016 28441 16028 28475
rect 16062 28472 16074 28475
rect 16666 28472 16672 28484
rect 16062 28444 16672 28472
rect 16062 28441 16074 28444
rect 16016 28435 16074 28441
rect 16666 28432 16672 28444
rect 16724 28432 16730 28484
rect 5258 28404 5264 28416
rect 5219 28376 5264 28404
rect 5258 28364 5264 28376
rect 5316 28364 5322 28416
rect 7374 28404 7380 28416
rect 7335 28376 7380 28404
rect 7374 28364 7380 28376
rect 7432 28364 7438 28416
rect 10226 28404 10232 28416
rect 10187 28376 10232 28404
rect 10226 28364 10232 28376
rect 10284 28364 10290 28416
rect 13449 28407 13507 28413
rect 13449 28373 13461 28407
rect 13495 28404 13507 28407
rect 13998 28404 14004 28416
rect 13495 28376 14004 28404
rect 13495 28373 13507 28376
rect 13449 28367 13507 28373
rect 13998 28364 14004 28376
rect 14056 28364 14062 28416
rect 1104 28314 18860 28336
rect 1104 28262 6880 28314
rect 6932 28262 6944 28314
rect 6996 28262 7008 28314
rect 7060 28262 7072 28314
rect 7124 28262 7136 28314
rect 7188 28262 12811 28314
rect 12863 28262 12875 28314
rect 12927 28262 12939 28314
rect 12991 28262 13003 28314
rect 13055 28262 13067 28314
rect 13119 28262 18860 28314
rect 1104 28240 18860 28262
rect 3786 28200 3792 28212
rect 3747 28172 3792 28200
rect 3786 28160 3792 28172
rect 3844 28160 3850 28212
rect 7177 28203 7235 28209
rect 7177 28169 7189 28203
rect 7223 28200 7235 28203
rect 7558 28200 7564 28212
rect 7223 28172 7564 28200
rect 7223 28169 7235 28172
rect 7177 28163 7235 28169
rect 7558 28160 7564 28172
rect 7616 28160 7622 28212
rect 7834 28200 7840 28212
rect 7795 28172 7840 28200
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 12526 28200 12532 28212
rect 12268 28172 12532 28200
rect 5258 28132 5264 28144
rect 4080 28104 5264 28132
rect 4080 28073 4108 28104
rect 5258 28092 5264 28104
rect 5316 28092 5322 28144
rect 7377 28135 7435 28141
rect 7377 28101 7389 28135
rect 7423 28101 7435 28135
rect 7377 28095 7435 28101
rect 4065 28067 4123 28073
rect 4065 28033 4077 28067
rect 4111 28033 4123 28067
rect 4065 28027 4123 28033
rect 4157 28067 4215 28073
rect 4157 28033 4169 28067
rect 4203 28033 4215 28067
rect 4157 28027 4215 28033
rect 4172 27996 4200 28027
rect 4246 28024 4252 28076
rect 4304 28064 4310 28076
rect 4304 28036 4349 28064
rect 4304 28024 4310 28036
rect 4430 28024 4436 28076
rect 4488 28064 4494 28076
rect 4798 28064 4804 28076
rect 4488 28036 4804 28064
rect 4488 28024 4494 28036
rect 4798 28024 4804 28036
rect 4856 28024 4862 28076
rect 7392 28064 7420 28095
rect 8113 28067 8171 28073
rect 8113 28064 8125 28067
rect 6886 28036 8125 28064
rect 4614 27996 4620 28008
rect 4172 27968 4620 27996
rect 4614 27956 4620 27968
rect 4672 27956 4678 28008
rect 6086 27956 6092 28008
rect 6144 27996 6150 28008
rect 6886 27996 6914 28036
rect 8113 28033 8125 28036
rect 8159 28064 8171 28067
rect 8294 28064 8300 28076
rect 8159 28036 8300 28064
rect 8159 28033 8171 28036
rect 8113 28027 8171 28033
rect 8294 28024 8300 28036
rect 8352 28024 8358 28076
rect 11882 28024 11888 28076
rect 11940 28064 11946 28076
rect 12268 28073 12296 28172
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 12710 28200 12716 28212
rect 12671 28172 12716 28200
rect 12710 28160 12716 28172
rect 12768 28160 12774 28212
rect 13173 28203 13231 28209
rect 13173 28169 13185 28203
rect 13219 28200 13231 28203
rect 13722 28200 13728 28212
rect 13219 28172 13728 28200
rect 13219 28169 13231 28172
rect 13173 28163 13231 28169
rect 13722 28160 13728 28172
rect 13780 28160 13786 28212
rect 16666 28200 16672 28212
rect 16627 28172 16672 28200
rect 16666 28160 16672 28172
rect 16724 28160 16730 28212
rect 13630 28132 13636 28144
rect 12360 28104 13636 28132
rect 12360 28073 12388 28104
rect 13630 28092 13636 28104
rect 13688 28092 13694 28144
rect 12069 28067 12127 28073
rect 12069 28064 12081 28067
rect 11940 28036 12081 28064
rect 11940 28024 11946 28036
rect 12069 28033 12081 28036
rect 12115 28033 12127 28067
rect 12069 28027 12127 28033
rect 12253 28067 12311 28073
rect 12253 28033 12265 28067
rect 12299 28033 12311 28067
rect 12253 28027 12311 28033
rect 12345 28067 12403 28073
rect 12345 28033 12357 28067
rect 12391 28033 12403 28067
rect 12345 28027 12403 28033
rect 12434 28024 12440 28076
rect 12492 28064 12498 28076
rect 14274 28064 14280 28076
rect 14332 28073 14338 28076
rect 12492 28036 12537 28064
rect 14244 28036 14280 28064
rect 12492 28024 12498 28036
rect 14274 28024 14280 28036
rect 14332 28027 14344 28073
rect 14553 28067 14611 28073
rect 14553 28033 14565 28067
rect 14599 28064 14611 28067
rect 15470 28064 15476 28076
rect 14599 28036 15476 28064
rect 14599 28033 14611 28036
rect 14553 28027 14611 28033
rect 14332 28024 14338 28027
rect 15470 28024 15476 28036
rect 15528 28024 15534 28076
rect 16850 28064 16856 28076
rect 16811 28036 16856 28064
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 6144 27968 6914 27996
rect 6144 27956 6150 27968
rect 7466 27956 7472 28008
rect 7524 27956 7530 28008
rect 7837 27999 7895 28005
rect 7837 27965 7849 27999
rect 7883 27996 7895 27999
rect 8202 27996 8208 28008
rect 7883 27968 8208 27996
rect 7883 27965 7895 27968
rect 7837 27959 7895 27965
rect 8202 27956 8208 27968
rect 8260 27996 8266 28008
rect 10410 27996 10416 28008
rect 8260 27968 10416 27996
rect 8260 27956 8266 27968
rect 10410 27956 10416 27968
rect 10468 27956 10474 28008
rect 7009 27931 7067 27937
rect 7009 27897 7021 27931
rect 7055 27928 7067 27931
rect 7484 27928 7512 27956
rect 7055 27900 7512 27928
rect 7055 27897 7067 27900
rect 7009 27891 7067 27897
rect 7193 27863 7251 27869
rect 7193 27829 7205 27863
rect 7239 27860 7251 27863
rect 7466 27860 7472 27872
rect 7239 27832 7472 27860
rect 7239 27829 7251 27832
rect 7193 27823 7251 27829
rect 7466 27820 7472 27832
rect 7524 27820 7530 27872
rect 8018 27860 8024 27872
rect 7979 27832 8024 27860
rect 8018 27820 8024 27832
rect 8076 27820 8082 27872
rect 1104 27770 18860 27792
rect 1104 27718 3915 27770
rect 3967 27718 3979 27770
rect 4031 27718 4043 27770
rect 4095 27718 4107 27770
rect 4159 27718 4171 27770
rect 4223 27718 9846 27770
rect 9898 27718 9910 27770
rect 9962 27718 9974 27770
rect 10026 27718 10038 27770
rect 10090 27718 10102 27770
rect 10154 27718 15776 27770
rect 15828 27718 15840 27770
rect 15892 27718 15904 27770
rect 15956 27718 15968 27770
rect 16020 27718 16032 27770
rect 16084 27718 18860 27770
rect 1104 27696 18860 27718
rect 5902 27656 5908 27668
rect 5863 27628 5908 27656
rect 5902 27616 5908 27628
rect 5960 27616 5966 27668
rect 8294 27656 8300 27668
rect 8255 27628 8300 27656
rect 8294 27616 8300 27628
rect 8352 27616 8358 27668
rect 13354 27656 13360 27668
rect 13315 27628 13360 27656
rect 13354 27616 13360 27628
rect 13412 27616 13418 27668
rect 14274 27656 14280 27668
rect 14235 27628 14280 27656
rect 14274 27616 14280 27628
rect 14332 27616 14338 27668
rect 9766 27548 9772 27600
rect 9824 27548 9830 27600
rect 10410 27548 10416 27600
rect 10468 27588 10474 27600
rect 10505 27591 10563 27597
rect 10505 27588 10517 27591
rect 10468 27560 10517 27588
rect 10468 27548 10474 27560
rect 10505 27557 10517 27560
rect 10551 27557 10563 27591
rect 13538 27588 13544 27600
rect 13499 27560 13544 27588
rect 10505 27551 10563 27557
rect 13538 27548 13544 27560
rect 13596 27548 13602 27600
rect 6917 27455 6975 27461
rect 6917 27421 6929 27455
rect 6963 27452 6975 27455
rect 9674 27452 9680 27464
rect 6963 27424 7328 27452
rect 9635 27424 9680 27452
rect 6963 27421 6975 27424
rect 6917 27415 6975 27421
rect 7300 27396 7328 27424
rect 9674 27412 9680 27424
rect 9732 27412 9738 27464
rect 9784 27461 9812 27548
rect 10226 27520 10232 27532
rect 9876 27492 10232 27520
rect 9876 27461 9904 27492
rect 10226 27480 10232 27492
rect 10284 27480 10290 27532
rect 9769 27455 9827 27461
rect 9769 27421 9781 27455
rect 9815 27421 9827 27455
rect 9769 27415 9827 27421
rect 9861 27455 9919 27461
rect 9861 27421 9873 27455
rect 9907 27421 9919 27455
rect 9861 27415 9919 27421
rect 10045 27455 10103 27461
rect 10045 27421 10057 27455
rect 10091 27452 10103 27455
rect 10318 27452 10324 27464
rect 10091 27424 10324 27452
rect 10091 27421 10103 27424
rect 10045 27415 10103 27421
rect 10318 27412 10324 27424
rect 10376 27412 10382 27464
rect 11330 27452 11336 27464
rect 11291 27424 11336 27452
rect 11330 27412 11336 27424
rect 11388 27412 11394 27464
rect 11606 27461 11612 27464
rect 11600 27452 11612 27461
rect 11519 27424 11612 27452
rect 11600 27415 11612 27424
rect 11664 27452 11670 27464
rect 12342 27452 12348 27464
rect 11664 27424 12348 27452
rect 11606 27412 11612 27415
rect 11664 27412 11670 27424
rect 12342 27412 12348 27424
rect 12400 27412 12406 27464
rect 13998 27412 14004 27464
rect 14056 27452 14062 27464
rect 14093 27455 14151 27461
rect 14093 27452 14105 27455
rect 14056 27424 14105 27452
rect 14056 27412 14062 27424
rect 14093 27421 14105 27424
rect 14139 27421 14151 27455
rect 14093 27415 14151 27421
rect 4430 27344 4436 27396
rect 4488 27384 4494 27396
rect 5537 27387 5595 27393
rect 5537 27384 5549 27387
rect 4488 27356 5549 27384
rect 4488 27344 4494 27356
rect 5537 27353 5549 27356
rect 5583 27353 5595 27387
rect 5718 27384 5724 27396
rect 5679 27356 5724 27384
rect 5537 27347 5595 27353
rect 5718 27344 5724 27356
rect 5776 27344 5782 27396
rect 7184 27387 7242 27393
rect 7184 27353 7196 27387
rect 7230 27353 7242 27387
rect 7184 27347 7242 27353
rect 4706 27276 4712 27328
rect 4764 27316 4770 27328
rect 5442 27316 5448 27328
rect 4764 27288 5448 27316
rect 4764 27276 4770 27288
rect 5442 27276 5448 27288
rect 5500 27276 5506 27328
rect 7208 27316 7236 27347
rect 7282 27344 7288 27396
rect 7340 27344 7346 27396
rect 10689 27387 10747 27393
rect 10689 27353 10701 27387
rect 10735 27384 10747 27387
rect 11882 27384 11888 27396
rect 10735 27356 11888 27384
rect 10735 27353 10747 27356
rect 10689 27347 10747 27353
rect 11882 27344 11888 27356
rect 11940 27344 11946 27396
rect 13173 27387 13231 27393
rect 13173 27384 13185 27387
rect 12728 27356 13185 27384
rect 7374 27316 7380 27328
rect 7208 27288 7380 27316
rect 7374 27276 7380 27288
rect 7432 27276 7438 27328
rect 9398 27316 9404 27328
rect 9359 27288 9404 27316
rect 9398 27276 9404 27288
rect 9456 27276 9462 27328
rect 12250 27276 12256 27328
rect 12308 27316 12314 27328
rect 12728 27325 12756 27356
rect 13173 27353 13185 27356
rect 13219 27353 13231 27387
rect 13173 27347 13231 27353
rect 13389 27387 13447 27393
rect 13389 27353 13401 27387
rect 13435 27384 13447 27387
rect 13814 27384 13820 27396
rect 13435 27356 13820 27384
rect 13435 27353 13447 27356
rect 13389 27347 13447 27353
rect 13814 27344 13820 27356
rect 13872 27344 13878 27396
rect 12713 27319 12771 27325
rect 12713 27316 12725 27319
rect 12308 27288 12725 27316
rect 12308 27276 12314 27288
rect 12713 27285 12725 27288
rect 12759 27285 12771 27319
rect 12713 27279 12771 27285
rect 1104 27226 18860 27248
rect 1104 27174 6880 27226
rect 6932 27174 6944 27226
rect 6996 27174 7008 27226
rect 7060 27174 7072 27226
rect 7124 27174 7136 27226
rect 7188 27174 12811 27226
rect 12863 27174 12875 27226
rect 12927 27174 12939 27226
rect 12991 27174 13003 27226
rect 13055 27174 13067 27226
rect 13119 27174 18860 27226
rect 1104 27152 18860 27174
rect 4706 27072 4712 27124
rect 4764 27112 4770 27124
rect 5077 27115 5135 27121
rect 5077 27112 5089 27115
rect 4764 27084 5089 27112
rect 4764 27072 4770 27084
rect 5077 27081 5089 27084
rect 5123 27112 5135 27115
rect 5718 27112 5724 27124
rect 5123 27084 5724 27112
rect 5123 27081 5135 27084
rect 5077 27075 5135 27081
rect 5718 27072 5724 27084
rect 5776 27072 5782 27124
rect 9674 27072 9680 27124
rect 9732 27112 9738 27124
rect 10505 27115 10563 27121
rect 10505 27112 10517 27115
rect 9732 27084 10517 27112
rect 9732 27072 9738 27084
rect 10505 27081 10517 27084
rect 10551 27081 10563 27115
rect 10505 27075 10563 27081
rect 11517 27115 11575 27121
rect 11517 27081 11529 27115
rect 11563 27112 11575 27115
rect 11606 27112 11612 27124
rect 11563 27084 11612 27112
rect 11563 27081 11575 27084
rect 11517 27075 11575 27081
rect 11606 27072 11612 27084
rect 11664 27072 11670 27124
rect 12161 27115 12219 27121
rect 12161 27081 12173 27115
rect 12207 27112 12219 27115
rect 12434 27112 12440 27124
rect 12207 27084 12440 27112
rect 12207 27081 12219 27084
rect 12161 27075 12219 27081
rect 12434 27072 12440 27084
rect 12492 27072 12498 27124
rect 16850 27072 16856 27124
rect 16908 27112 16914 27124
rect 17037 27115 17095 27121
rect 17037 27112 17049 27115
rect 16908 27084 17049 27112
rect 16908 27072 16914 27084
rect 17037 27081 17049 27084
rect 17083 27081 17095 27115
rect 17037 27075 17095 27081
rect 7282 27004 7288 27056
rect 7340 27044 7346 27056
rect 9398 27053 9404 27056
rect 9392 27044 9404 27053
rect 7340 27016 8708 27044
rect 9359 27016 9404 27044
rect 7340 27004 7346 27016
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 4522 26976 4528 26988
rect 1719 26948 4528 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 4522 26936 4528 26948
rect 4580 26936 4586 26988
rect 4982 26976 4988 26988
rect 4943 26948 4988 26976
rect 4982 26936 4988 26948
rect 5040 26936 5046 26988
rect 8386 26976 8392 26988
rect 8444 26985 8450 26988
rect 8680 26985 8708 27016
rect 9392 27007 9404 27016
rect 9398 27004 9404 27007
rect 9456 27004 9462 27056
rect 12526 27004 12532 27056
rect 12584 27044 12590 27056
rect 12621 27047 12679 27053
rect 12621 27044 12633 27047
rect 12584 27016 12633 27044
rect 12584 27004 12590 27016
rect 12621 27013 12633 27016
rect 12667 27044 12679 27047
rect 13354 27044 13360 27056
rect 12667 27016 13360 27044
rect 12667 27013 12679 27016
rect 12621 27007 12679 27013
rect 13354 27004 13360 27016
rect 13412 27004 13418 27056
rect 8356 26948 8392 26976
rect 8386 26936 8392 26948
rect 8444 26939 8456 26985
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26976 8723 26979
rect 9125 26979 9183 26985
rect 9125 26976 9137 26979
rect 8711 26948 9137 26976
rect 8711 26945 8723 26948
rect 8665 26939 8723 26945
rect 9125 26945 9137 26948
rect 9171 26976 9183 26979
rect 9766 26976 9772 26988
rect 9171 26948 9772 26976
rect 9171 26945 9183 26948
rect 9125 26939 9183 26945
rect 8444 26936 8450 26939
rect 9766 26936 9772 26948
rect 9824 26936 9830 26988
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26976 11759 26979
rect 12066 26976 12072 26988
rect 11747 26948 12072 26976
rect 11747 26945 11759 26948
rect 11701 26939 11759 26945
rect 12066 26936 12072 26948
rect 12124 26936 12130 26988
rect 12250 26936 12256 26988
rect 12308 26976 12314 26988
rect 12345 26979 12403 26985
rect 12345 26976 12357 26979
rect 12308 26948 12357 26976
rect 12308 26936 12314 26948
rect 12345 26945 12357 26948
rect 12391 26945 12403 26979
rect 16758 26976 16764 26988
rect 16719 26948 16764 26976
rect 12345 26939 12403 26945
rect 16758 26936 16764 26948
rect 16816 26936 16822 26988
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26976 16911 26979
rect 16942 26976 16948 26988
rect 16899 26948 16948 26976
rect 16899 26945 16911 26948
rect 16853 26939 16911 26945
rect 16942 26936 16948 26948
rect 17000 26936 17006 26988
rect 12529 26911 12587 26917
rect 12529 26877 12541 26911
rect 12575 26908 12587 26911
rect 12618 26908 12624 26920
rect 12575 26880 12624 26908
rect 12575 26877 12587 26880
rect 12529 26871 12587 26877
rect 12618 26868 12624 26880
rect 12676 26868 12682 26920
rect 7285 26843 7343 26849
rect 7285 26840 7297 26843
rect 6886 26812 7297 26840
rect 1486 26772 1492 26784
rect 1447 26744 1492 26772
rect 1486 26732 1492 26744
rect 1544 26732 1550 26784
rect 4430 26732 4436 26784
rect 4488 26772 4494 26784
rect 6886 26772 6914 26812
rect 7285 26809 7297 26812
rect 7331 26840 7343 26843
rect 7466 26840 7472 26852
rect 7331 26812 7472 26840
rect 7331 26809 7343 26812
rect 7285 26803 7343 26809
rect 7466 26800 7472 26812
rect 7524 26800 7530 26852
rect 11698 26800 11704 26852
rect 11756 26840 11762 26852
rect 13446 26840 13452 26852
rect 11756 26812 13452 26840
rect 11756 26800 11762 26812
rect 13446 26800 13452 26812
rect 13504 26800 13510 26852
rect 4488 26744 6914 26772
rect 4488 26732 4494 26744
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 12492 26744 12537 26772
rect 12492 26732 12498 26744
rect 1104 26682 18860 26704
rect 1104 26630 3915 26682
rect 3967 26630 3979 26682
rect 4031 26630 4043 26682
rect 4095 26630 4107 26682
rect 4159 26630 4171 26682
rect 4223 26630 9846 26682
rect 9898 26630 9910 26682
rect 9962 26630 9974 26682
rect 10026 26630 10038 26682
rect 10090 26630 10102 26682
rect 10154 26630 15776 26682
rect 15828 26630 15840 26682
rect 15892 26630 15904 26682
rect 15956 26630 15968 26682
rect 16020 26630 16032 26682
rect 16084 26630 18860 26682
rect 1104 26608 18860 26630
rect 4433 26571 4491 26577
rect 4433 26537 4445 26571
rect 4479 26568 4491 26571
rect 5534 26568 5540 26580
rect 4479 26540 5540 26568
rect 4479 26537 4491 26540
rect 4433 26531 4491 26537
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 7745 26571 7803 26577
rect 5644 26540 7696 26568
rect 1670 26460 1676 26512
rect 1728 26500 1734 26512
rect 5644 26500 5672 26540
rect 1728 26472 5672 26500
rect 7668 26500 7696 26540
rect 7745 26537 7757 26571
rect 7791 26568 7803 26571
rect 8018 26568 8024 26580
rect 7791 26540 8024 26568
rect 7791 26537 7803 26540
rect 7745 26531 7803 26537
rect 8018 26528 8024 26540
rect 8076 26528 8082 26580
rect 8386 26568 8392 26580
rect 8347 26540 8392 26568
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 12066 26568 12072 26580
rect 12027 26540 12072 26568
rect 12066 26528 12072 26540
rect 12124 26528 12130 26580
rect 11241 26503 11299 26509
rect 7668 26472 9260 26500
rect 1728 26460 1734 26472
rect 3602 26392 3608 26444
rect 3660 26432 3666 26444
rect 7282 26432 7288 26444
rect 3660 26404 5948 26432
rect 3660 26392 3666 26404
rect 4430 26324 4436 26376
rect 4488 26364 4494 26376
rect 4571 26367 4629 26373
rect 4571 26364 4583 26367
rect 4488 26336 4583 26364
rect 4488 26324 4494 26336
rect 4571 26333 4583 26336
rect 4617 26333 4629 26367
rect 4571 26327 4629 26333
rect 4706 26324 4712 26376
rect 4764 26364 4770 26376
rect 4984 26367 5042 26373
rect 4764 26336 4809 26364
rect 4764 26324 4770 26336
rect 4984 26333 4996 26367
rect 5030 26333 5042 26367
rect 4984 26327 5042 26333
rect 4801 26299 4859 26305
rect 4801 26265 4813 26299
rect 4847 26265 4859 26299
rect 5000 26296 5028 26327
rect 5074 26324 5080 26376
rect 5132 26364 5138 26376
rect 5920 26364 5948 26404
rect 7208 26404 7288 26432
rect 6917 26367 6975 26373
rect 6917 26364 6929 26367
rect 5132 26336 5177 26364
rect 5920 26336 6929 26364
rect 5132 26324 5138 26336
rect 6917 26333 6929 26336
rect 6963 26364 6975 26367
rect 7208 26364 7236 26404
rect 7282 26392 7288 26404
rect 7340 26392 7346 26444
rect 7374 26364 7380 26376
rect 6963 26336 7236 26364
rect 7335 26336 7380 26364
rect 6963 26333 6975 26336
rect 6917 26327 6975 26333
rect 7374 26324 7380 26336
rect 7432 26324 7438 26376
rect 7558 26364 7564 26376
rect 7519 26336 7564 26364
rect 7558 26324 7564 26336
rect 7616 26324 7622 26376
rect 8018 26324 8024 26376
rect 8076 26364 8082 26376
rect 8205 26367 8263 26373
rect 8205 26364 8217 26367
rect 8076 26336 8217 26364
rect 8076 26324 8082 26336
rect 8205 26333 8217 26336
rect 8251 26333 8263 26367
rect 8386 26364 8392 26376
rect 8347 26336 8392 26364
rect 8205 26327 8263 26333
rect 8386 26324 8392 26336
rect 8444 26324 8450 26376
rect 9232 26373 9260 26472
rect 11241 26469 11253 26503
rect 11287 26469 11299 26503
rect 11241 26463 11299 26469
rect 9766 26392 9772 26444
rect 9824 26432 9830 26444
rect 9861 26435 9919 26441
rect 9861 26432 9873 26435
rect 9824 26404 9873 26432
rect 9824 26392 9830 26404
rect 9861 26401 9873 26404
rect 9907 26401 9919 26435
rect 11256 26432 11284 26463
rect 12434 26432 12440 26444
rect 11256 26404 12440 26432
rect 9861 26395 9919 26401
rect 12434 26392 12440 26404
rect 12492 26432 12498 26444
rect 12492 26404 12537 26432
rect 12492 26392 12498 26404
rect 9125 26367 9183 26373
rect 9125 26333 9137 26367
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 11698 26364 11704 26376
rect 9217 26327 9275 26333
rect 9324 26336 11704 26364
rect 5166 26296 5172 26308
rect 5000 26268 5172 26296
rect 4801 26259 4859 26265
rect 4816 26228 4844 26259
rect 5166 26256 5172 26268
rect 5224 26256 5230 26308
rect 6362 26256 6368 26308
rect 6420 26296 6426 26308
rect 6650 26299 6708 26305
rect 6650 26296 6662 26299
rect 6420 26268 6662 26296
rect 6420 26256 6426 26268
rect 6650 26265 6662 26268
rect 6696 26265 6708 26299
rect 9140 26296 9168 26327
rect 9324 26296 9352 26336
rect 11698 26324 11704 26336
rect 11756 26324 11762 26376
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26364 12311 26367
rect 14090 26364 14096 26376
rect 12299 26336 14096 26364
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 14090 26324 14096 26336
rect 14148 26324 14154 26376
rect 9140 26268 9352 26296
rect 9401 26299 9459 26305
rect 6650 26259 6708 26265
rect 9401 26265 9413 26299
rect 9447 26296 9459 26299
rect 10128 26299 10186 26305
rect 9447 26268 9674 26296
rect 9447 26265 9459 26268
rect 9401 26259 9459 26265
rect 5350 26228 5356 26240
rect 4816 26200 5356 26228
rect 5350 26188 5356 26200
rect 5408 26228 5414 26240
rect 5537 26231 5595 26237
rect 5537 26228 5549 26231
rect 5408 26200 5549 26228
rect 5408 26188 5414 26200
rect 5537 26197 5549 26200
rect 5583 26197 5595 26231
rect 9646 26228 9674 26268
rect 10128 26265 10140 26299
rect 10174 26296 10186 26299
rect 10410 26296 10416 26308
rect 10174 26268 10416 26296
rect 10174 26265 10186 26268
rect 10128 26259 10186 26265
rect 10410 26256 10416 26268
rect 10468 26256 10474 26308
rect 10686 26228 10692 26240
rect 9646 26200 10692 26228
rect 5537 26191 5595 26197
rect 10686 26188 10692 26200
rect 10744 26188 10750 26240
rect 1104 26138 18860 26160
rect 1104 26086 6880 26138
rect 6932 26086 6944 26138
rect 6996 26086 7008 26138
rect 7060 26086 7072 26138
rect 7124 26086 7136 26138
rect 7188 26086 12811 26138
rect 12863 26086 12875 26138
rect 12927 26086 12939 26138
rect 12991 26086 13003 26138
rect 13055 26086 13067 26138
rect 13119 26086 18860 26138
rect 1104 26064 18860 26086
rect 6362 26024 6368 26036
rect 6323 25996 6368 26024
rect 6362 25984 6368 25996
rect 6420 25984 6426 26036
rect 8021 26027 8079 26033
rect 8021 25993 8033 26027
rect 8067 26024 8079 26027
rect 8386 26024 8392 26036
rect 8067 25996 8392 26024
rect 8067 25993 8079 25996
rect 8021 25987 8079 25993
rect 8386 25984 8392 25996
rect 8444 25984 8450 26036
rect 9861 26027 9919 26033
rect 9861 25993 9873 26027
rect 9907 26024 9919 26027
rect 10318 26024 10324 26036
rect 9907 25996 10324 26024
rect 9907 25993 9919 25996
rect 9861 25987 9919 25993
rect 10318 25984 10324 25996
rect 10376 25984 10382 26036
rect 10410 25984 10416 26036
rect 10468 26024 10474 26036
rect 10505 26027 10563 26033
rect 10505 26024 10517 26027
rect 10468 25996 10517 26024
rect 10468 25984 10474 25996
rect 10505 25993 10517 25996
rect 10551 25993 10563 26027
rect 10505 25987 10563 25993
rect 11517 26027 11575 26033
rect 11517 25993 11529 26027
rect 11563 26024 11575 26027
rect 12618 26024 12624 26036
rect 11563 25996 12624 26024
rect 11563 25993 11575 25996
rect 11517 25987 11575 25993
rect 12618 25984 12624 25996
rect 12676 25984 12682 26036
rect 5626 25916 5632 25968
rect 5684 25956 5690 25968
rect 6641 25959 6699 25965
rect 6641 25956 6653 25959
rect 5684 25928 6653 25956
rect 5684 25916 5690 25928
rect 6641 25925 6653 25928
rect 6687 25956 6699 25959
rect 7282 25956 7288 25968
rect 6687 25928 7288 25956
rect 6687 25925 6699 25928
rect 6641 25919 6699 25925
rect 7282 25916 7288 25928
rect 7340 25916 7346 25968
rect 11330 25916 11336 25968
rect 11388 25956 11394 25968
rect 11388 25928 12940 25956
rect 11388 25916 11394 25928
rect 3602 25888 3608 25900
rect 3563 25860 3608 25888
rect 3602 25848 3608 25860
rect 3660 25848 3666 25900
rect 3694 25848 3700 25900
rect 3752 25888 3758 25900
rect 3861 25891 3919 25897
rect 3861 25888 3873 25891
rect 3752 25860 3873 25888
rect 3752 25848 3758 25860
rect 3861 25857 3873 25860
rect 3907 25857 3919 25891
rect 3861 25851 3919 25857
rect 6365 25891 6423 25897
rect 6365 25857 6377 25891
rect 6411 25888 6423 25891
rect 6411 25860 6914 25888
rect 6411 25857 6423 25860
rect 6365 25851 6423 25857
rect 6886 25832 6914 25860
rect 7374 25848 7380 25900
rect 7432 25888 7438 25900
rect 7745 25891 7803 25897
rect 7745 25888 7757 25891
rect 7432 25860 7757 25888
rect 7432 25848 7438 25860
rect 7745 25857 7757 25860
rect 7791 25857 7803 25891
rect 7745 25851 7803 25857
rect 9953 25891 10011 25897
rect 9953 25857 9965 25891
rect 9999 25888 10011 25891
rect 10410 25888 10416 25900
rect 9999 25860 10416 25888
rect 9999 25857 10011 25860
rect 9953 25851 10011 25857
rect 10410 25848 10416 25860
rect 10468 25848 10474 25900
rect 10686 25888 10692 25900
rect 10647 25860 10692 25888
rect 10686 25848 10692 25860
rect 10744 25848 10750 25900
rect 12641 25891 12699 25897
rect 12641 25857 12653 25891
rect 12687 25888 12699 25891
rect 12802 25888 12808 25900
rect 12687 25860 12808 25888
rect 12687 25857 12699 25860
rect 12641 25851 12699 25857
rect 12802 25848 12808 25860
rect 12860 25848 12866 25900
rect 12912 25897 12940 25928
rect 12897 25891 12955 25897
rect 12897 25857 12909 25891
rect 12943 25857 12955 25891
rect 15470 25888 15476 25900
rect 15431 25860 15476 25888
rect 12897 25851 12955 25857
rect 15470 25848 15476 25860
rect 15528 25848 15534 25900
rect 16574 25848 16580 25900
rect 16632 25888 16638 25900
rect 16669 25891 16727 25897
rect 16669 25888 16681 25891
rect 16632 25860 16681 25888
rect 16632 25848 16638 25860
rect 16669 25857 16681 25860
rect 16715 25857 16727 25891
rect 16669 25851 16727 25857
rect 6886 25792 6920 25832
rect 6914 25780 6920 25792
rect 6972 25820 6978 25832
rect 7558 25820 7564 25832
rect 6972 25792 7564 25820
rect 6972 25780 6978 25792
rect 7558 25780 7564 25792
rect 7616 25820 7622 25832
rect 7837 25823 7895 25829
rect 7837 25820 7849 25823
rect 7616 25792 7849 25820
rect 7616 25780 7622 25792
rect 7837 25789 7849 25792
rect 7883 25789 7895 25823
rect 7837 25783 7895 25789
rect 8021 25823 8079 25829
rect 8021 25789 8033 25823
rect 8067 25820 8079 25823
rect 11606 25820 11612 25832
rect 8067 25792 11612 25820
rect 8067 25789 8079 25792
rect 8021 25783 8079 25789
rect 11606 25780 11612 25792
rect 11664 25780 11670 25832
rect 16758 25820 16764 25832
rect 16719 25792 16764 25820
rect 16758 25780 16764 25792
rect 16816 25780 16822 25832
rect 5258 25712 5264 25764
rect 5316 25752 5322 25764
rect 6457 25755 6515 25761
rect 6457 25752 6469 25755
rect 5316 25724 6469 25752
rect 5316 25712 5322 25724
rect 6457 25721 6469 25724
rect 6503 25721 6515 25755
rect 17954 25752 17960 25764
rect 6457 25715 6515 25721
rect 16868 25724 17960 25752
rect 4982 25684 4988 25696
rect 4943 25656 4988 25684
rect 4982 25644 4988 25656
rect 5040 25644 5046 25696
rect 15562 25644 15568 25696
rect 15620 25684 15626 25696
rect 16868 25693 16896 25724
rect 17954 25712 17960 25724
rect 18012 25712 18018 25764
rect 15657 25687 15715 25693
rect 15657 25684 15669 25687
rect 15620 25656 15669 25684
rect 15620 25644 15626 25656
rect 15657 25653 15669 25656
rect 15703 25653 15715 25687
rect 15657 25647 15715 25653
rect 16853 25687 16911 25693
rect 16853 25653 16865 25687
rect 16899 25653 16911 25687
rect 17034 25684 17040 25696
rect 16995 25656 17040 25684
rect 16853 25647 16911 25653
rect 17034 25644 17040 25656
rect 17092 25644 17098 25696
rect 1104 25594 18860 25616
rect 1104 25542 3915 25594
rect 3967 25542 3979 25594
rect 4031 25542 4043 25594
rect 4095 25542 4107 25594
rect 4159 25542 4171 25594
rect 4223 25542 9846 25594
rect 9898 25542 9910 25594
rect 9962 25542 9974 25594
rect 10026 25542 10038 25594
rect 10090 25542 10102 25594
rect 10154 25542 15776 25594
rect 15828 25542 15840 25594
rect 15892 25542 15904 25594
rect 15956 25542 15968 25594
rect 16020 25542 16032 25594
rect 16084 25542 18860 25594
rect 1104 25520 18860 25542
rect 3694 25440 3700 25492
rect 3752 25480 3758 25492
rect 3789 25483 3847 25489
rect 3789 25480 3801 25483
rect 3752 25452 3801 25480
rect 3752 25440 3758 25452
rect 3789 25449 3801 25452
rect 3835 25449 3847 25483
rect 5258 25480 5264 25492
rect 5219 25452 5264 25480
rect 3789 25443 3847 25449
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 5626 25440 5632 25492
rect 5684 25480 5690 25492
rect 6181 25483 6239 25489
rect 6181 25480 6193 25483
rect 5684 25452 6193 25480
rect 5684 25440 5690 25452
rect 6181 25449 6193 25452
rect 6227 25449 6239 25483
rect 6181 25443 6239 25449
rect 6365 25483 6423 25489
rect 6365 25449 6377 25483
rect 6411 25480 6423 25483
rect 6914 25480 6920 25492
rect 6411 25452 6920 25480
rect 6411 25449 6423 25452
rect 6365 25443 6423 25449
rect 6914 25440 6920 25452
rect 6972 25440 6978 25492
rect 12802 25440 12808 25492
rect 12860 25480 12866 25492
rect 13265 25483 13323 25489
rect 13265 25480 13277 25483
rect 12860 25452 13277 25480
rect 12860 25440 12866 25452
rect 13265 25449 13277 25452
rect 13311 25449 13323 25483
rect 13265 25443 13323 25449
rect 16577 25483 16635 25489
rect 16577 25449 16589 25483
rect 16623 25480 16635 25483
rect 16666 25480 16672 25492
rect 16623 25452 16672 25480
rect 16623 25449 16635 25452
rect 16577 25443 16635 25449
rect 16666 25440 16672 25452
rect 16724 25480 16730 25492
rect 16850 25480 16856 25492
rect 16724 25452 16856 25480
rect 16724 25440 16730 25452
rect 16850 25440 16856 25452
rect 16908 25440 16914 25492
rect 3234 25372 3240 25424
rect 3292 25412 3298 25424
rect 3292 25384 9812 25412
rect 3292 25372 3298 25384
rect 4982 25344 4988 25356
rect 4080 25316 4988 25344
rect 3694 25236 3700 25288
rect 3752 25276 3758 25288
rect 4080 25285 4108 25316
rect 4982 25304 4988 25316
rect 5040 25304 5046 25356
rect 4065 25279 4123 25285
rect 4065 25276 4077 25279
rect 3752 25248 4077 25276
rect 3752 25236 3758 25248
rect 4065 25245 4077 25248
rect 4111 25245 4123 25279
rect 4065 25239 4123 25245
rect 4157 25279 4215 25285
rect 4157 25245 4169 25279
rect 4203 25245 4215 25279
rect 4157 25239 4215 25245
rect 4172 25208 4200 25239
rect 4246 25236 4252 25288
rect 4304 25276 4310 25288
rect 4433 25279 4491 25285
rect 4304 25248 4349 25276
rect 4304 25236 4310 25248
rect 4433 25245 4445 25279
rect 4479 25276 4491 25279
rect 4798 25276 4804 25288
rect 4479 25248 4804 25276
rect 4479 25245 4491 25248
rect 4433 25239 4491 25245
rect 4798 25236 4804 25248
rect 4856 25236 4862 25288
rect 5261 25279 5319 25285
rect 5261 25245 5273 25279
rect 5307 25276 5319 25279
rect 5350 25276 5356 25288
rect 5307 25248 5356 25276
rect 5307 25245 5319 25248
rect 5261 25239 5319 25245
rect 5350 25236 5356 25248
rect 5408 25236 5414 25288
rect 5537 25279 5595 25285
rect 5537 25245 5549 25279
rect 5583 25276 5595 25279
rect 5718 25276 5724 25288
rect 5583 25248 5724 25276
rect 5583 25245 5595 25248
rect 5537 25239 5595 25245
rect 5718 25236 5724 25248
rect 5776 25276 5782 25288
rect 9784 25285 9812 25384
rect 11606 25372 11612 25424
rect 11664 25412 11670 25424
rect 12066 25412 12072 25424
rect 11664 25384 12072 25412
rect 11664 25372 11670 25384
rect 12066 25372 12072 25384
rect 12124 25412 12130 25424
rect 16298 25412 16304 25424
rect 12124 25384 16304 25412
rect 12124 25372 12130 25384
rect 16298 25372 16304 25384
rect 16356 25372 16362 25424
rect 11977 25347 12035 25353
rect 11977 25313 11989 25347
rect 12023 25344 12035 25347
rect 12250 25344 12256 25356
rect 12023 25316 12256 25344
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 12250 25304 12256 25316
rect 12308 25304 12314 25356
rect 16574 25344 16580 25356
rect 15697 25316 16580 25344
rect 9677 25279 9735 25285
rect 5776 25248 6132 25276
rect 5776 25236 5782 25248
rect 4614 25208 4620 25220
rect 4172 25180 4620 25208
rect 4614 25168 4620 25180
rect 4672 25168 4678 25220
rect 5368 25208 5396 25236
rect 5997 25211 6055 25217
rect 5997 25208 6009 25211
rect 5368 25180 6009 25208
rect 5997 25177 6009 25180
rect 6043 25177 6055 25211
rect 6104 25208 6132 25248
rect 9677 25245 9689 25279
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 9769 25279 9827 25285
rect 9769 25245 9781 25279
rect 9815 25245 9827 25279
rect 9769 25239 9827 25245
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25276 11023 25279
rect 11609 25279 11667 25285
rect 11609 25276 11621 25279
rect 11011 25248 11621 25276
rect 11011 25245 11023 25248
rect 10965 25239 11023 25245
rect 11609 25245 11621 25248
rect 11655 25245 11667 25279
rect 11609 25239 11667 25245
rect 6197 25211 6255 25217
rect 6197 25208 6209 25211
rect 6104 25180 6209 25208
rect 5997 25171 6055 25177
rect 6197 25177 6209 25180
rect 6243 25177 6255 25211
rect 9692 25208 9720 25239
rect 11790 25236 11796 25288
rect 11848 25276 11854 25288
rect 12526 25276 12532 25288
rect 11848 25248 11941 25276
rect 12487 25248 12532 25276
rect 11848 25236 11854 25248
rect 12526 25236 12532 25248
rect 12584 25236 12590 25288
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25245 12679 25279
rect 12621 25239 12679 25245
rect 12805 25279 12863 25285
rect 12805 25245 12817 25279
rect 12851 25276 12863 25279
rect 13449 25279 13507 25285
rect 13449 25276 13461 25279
rect 12851 25248 13461 25276
rect 12851 25245 12863 25248
rect 12805 25239 12863 25245
rect 13449 25245 13461 25248
rect 13495 25245 13507 25279
rect 14458 25276 14464 25288
rect 14419 25248 14464 25276
rect 13449 25239 13507 25245
rect 9953 25211 10011 25217
rect 9692 25180 9812 25208
rect 6197 25171 6255 25177
rect 5445 25143 5503 25149
rect 5445 25109 5457 25143
rect 5491 25140 5503 25143
rect 5626 25140 5632 25152
rect 5491 25112 5632 25140
rect 5491 25109 5503 25112
rect 5445 25103 5503 25109
rect 5626 25100 5632 25112
rect 5684 25100 5690 25152
rect 9784 25140 9812 25180
rect 9953 25177 9965 25211
rect 9999 25208 10011 25211
rect 11514 25208 11520 25220
rect 9999 25180 11520 25208
rect 9999 25177 10011 25180
rect 9953 25171 10011 25177
rect 11514 25168 11520 25180
rect 11572 25168 11578 25220
rect 11808 25208 11836 25236
rect 12636 25208 12664 25239
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 11808 25180 12664 25208
rect 10410 25140 10416 25152
rect 9784 25112 10416 25140
rect 10410 25100 10416 25112
rect 10468 25100 10474 25152
rect 11146 25140 11152 25152
rect 11107 25112 11152 25140
rect 11146 25100 11152 25112
rect 11204 25100 11210 25152
rect 11330 25100 11336 25152
rect 11388 25140 11394 25152
rect 11808 25140 11836 25180
rect 11388 25112 11836 25140
rect 14645 25143 14703 25149
rect 11388 25100 11394 25112
rect 14645 25109 14657 25143
rect 14691 25140 14703 25143
rect 14826 25140 14832 25152
rect 14691 25112 14832 25140
rect 14691 25109 14703 25112
rect 14645 25103 14703 25109
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 15286 25140 15292 25152
rect 15247 25112 15292 25140
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 15488 25140 15516 25239
rect 15562 25236 15568 25288
rect 15620 25276 15626 25288
rect 15620 25248 15665 25276
rect 15620 25236 15626 25248
rect 15697 25217 15725 25316
rect 16574 25304 16580 25316
rect 16632 25304 16638 25356
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25276 15991 25279
rect 16666 25276 16672 25288
rect 15979 25248 16672 25276
rect 15979 25245 15991 25248
rect 15933 25239 15991 25245
rect 16666 25236 16672 25248
rect 16724 25236 16730 25288
rect 15657 25211 15725 25217
rect 15657 25177 15669 25211
rect 15703 25180 15725 25211
rect 15795 25211 15853 25217
rect 15703 25177 15715 25180
rect 15657 25171 15715 25177
rect 15795 25177 15807 25211
rect 15841 25208 15853 25211
rect 16298 25208 16304 25220
rect 15841 25180 16304 25208
rect 15841 25177 15853 25180
rect 15795 25171 15853 25177
rect 16298 25168 16304 25180
rect 16356 25168 16362 25220
rect 16758 25208 16764 25220
rect 16719 25180 16764 25208
rect 16758 25168 16764 25180
rect 16816 25168 16822 25220
rect 16393 25143 16451 25149
rect 16393 25140 16405 25143
rect 15488 25112 16405 25140
rect 16393 25109 16405 25112
rect 16439 25109 16451 25143
rect 16393 25103 16451 25109
rect 16561 25143 16619 25149
rect 16561 25109 16573 25143
rect 16607 25140 16619 25143
rect 17126 25140 17132 25152
rect 16607 25112 17132 25140
rect 16607 25109 16619 25112
rect 16561 25103 16619 25109
rect 17126 25100 17132 25112
rect 17184 25100 17190 25152
rect 1104 25050 18860 25072
rect 1104 24998 6880 25050
rect 6932 24998 6944 25050
rect 6996 24998 7008 25050
rect 7060 24998 7072 25050
rect 7124 24998 7136 25050
rect 7188 24998 12811 25050
rect 12863 24998 12875 25050
rect 12927 24998 12939 25050
rect 12991 24998 13003 25050
rect 13055 24998 13067 25050
rect 13119 24998 18860 25050
rect 1104 24976 18860 24998
rect 12526 24896 12532 24948
rect 12584 24936 12590 24948
rect 12897 24939 12955 24945
rect 12897 24936 12909 24939
rect 12584 24908 12909 24936
rect 12584 24896 12590 24908
rect 12897 24905 12909 24908
rect 12943 24905 12955 24939
rect 12897 24899 12955 24905
rect 14277 24939 14335 24945
rect 14277 24905 14289 24939
rect 14323 24936 14335 24939
rect 14458 24936 14464 24948
rect 14323 24908 14464 24936
rect 14323 24905 14335 24908
rect 14277 24899 14335 24905
rect 14458 24896 14464 24908
rect 14516 24896 14522 24948
rect 16942 24936 16948 24948
rect 14568 24908 16948 24936
rect 11146 24828 11152 24880
rect 11204 24868 11210 24880
rect 11762 24871 11820 24877
rect 11762 24868 11774 24871
rect 11204 24840 11774 24868
rect 11204 24828 11210 24840
rect 11762 24837 11774 24840
rect 11808 24837 11820 24871
rect 11762 24831 11820 24837
rect 5074 24800 5080 24812
rect 5035 24772 5080 24800
rect 5074 24760 5080 24772
rect 5132 24760 5138 24812
rect 5166 24760 5172 24812
rect 5224 24800 5230 24812
rect 5261 24803 5319 24809
rect 5261 24800 5273 24803
rect 5224 24772 5273 24800
rect 5224 24760 5230 24772
rect 5261 24769 5273 24772
rect 5307 24769 5319 24803
rect 5261 24763 5319 24769
rect 5350 24760 5356 24812
rect 5408 24800 5414 24812
rect 5445 24803 5503 24809
rect 5445 24800 5457 24803
rect 5408 24772 5457 24800
rect 5408 24760 5414 24772
rect 5445 24769 5457 24772
rect 5491 24769 5503 24803
rect 5626 24800 5632 24812
rect 5587 24772 5632 24800
rect 5445 24763 5503 24769
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 5810 24800 5816 24812
rect 5771 24772 5816 24800
rect 5810 24760 5816 24772
rect 5868 24760 5874 24812
rect 14093 24803 14151 24809
rect 14093 24769 14105 24803
rect 14139 24800 14151 24803
rect 14568 24800 14596 24908
rect 16942 24896 16948 24908
rect 17000 24896 17006 24948
rect 14936 24840 15424 24868
rect 14936 24800 14964 24840
rect 14139 24772 14596 24800
rect 14660 24772 14964 24800
rect 15004 24803 15062 24809
rect 14139 24769 14151 24772
rect 14093 24763 14151 24769
rect 14660 24744 14688 24772
rect 15004 24769 15016 24803
rect 15050 24800 15062 24803
rect 15286 24800 15292 24812
rect 15050 24772 15292 24800
rect 15050 24769 15062 24772
rect 15004 24763 15062 24769
rect 15286 24760 15292 24772
rect 15344 24760 15350 24812
rect 15396 24800 15424 24840
rect 16666 24800 16672 24812
rect 15396 24772 16160 24800
rect 16627 24772 16672 24800
rect 5534 24692 5540 24744
rect 5592 24732 5598 24744
rect 11517 24735 11575 24741
rect 5592 24704 5637 24732
rect 5592 24692 5598 24704
rect 11517 24701 11529 24735
rect 11563 24701 11575 24735
rect 11517 24695 11575 24701
rect 13909 24735 13967 24741
rect 13909 24701 13921 24735
rect 13955 24732 13967 24735
rect 14642 24732 14648 24744
rect 13955 24704 14648 24732
rect 13955 24701 13967 24704
rect 13909 24695 13967 24701
rect 11532 24596 11560 24695
rect 14642 24692 14648 24704
rect 14700 24692 14706 24744
rect 14737 24735 14795 24741
rect 14737 24701 14749 24735
rect 14783 24701 14795 24735
rect 14737 24695 14795 24701
rect 16132 24732 16160 24772
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 16850 24800 16856 24812
rect 16811 24772 16856 24800
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 16945 24803 17003 24809
rect 16945 24769 16957 24803
rect 16991 24800 17003 24803
rect 17034 24800 17040 24812
rect 16991 24772 17040 24800
rect 16991 24769 17003 24772
rect 16945 24763 17003 24769
rect 17034 24760 17040 24772
rect 17092 24760 17098 24812
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24769 17187 24803
rect 17129 24763 17187 24769
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24800 17923 24803
rect 18046 24800 18052 24812
rect 17911 24772 18052 24800
rect 17911 24769 17923 24772
rect 17865 24763 17923 24769
rect 17144 24732 17172 24763
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 18196 24772 18241 24800
rect 18196 24760 18202 24772
rect 16132 24704 17172 24732
rect 12250 24596 12256 24608
rect 11532 24568 12256 24596
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 14752 24596 14780 24695
rect 16132 24673 16160 24704
rect 17402 24692 17408 24744
rect 17460 24732 17466 24744
rect 17957 24735 18015 24741
rect 17957 24732 17969 24735
rect 17460 24704 17969 24732
rect 17460 24692 17466 24704
rect 17957 24701 17969 24704
rect 18003 24701 18015 24735
rect 17957 24695 18015 24701
rect 16117 24667 16175 24673
rect 16117 24633 16129 24667
rect 16163 24633 16175 24667
rect 16117 24627 16175 24633
rect 17037 24667 17095 24673
rect 17037 24633 17049 24667
rect 17083 24664 17095 24667
rect 17681 24667 17739 24673
rect 17681 24664 17693 24667
rect 17083 24636 17693 24664
rect 17083 24633 17095 24636
rect 17037 24627 17095 24633
rect 17681 24633 17693 24636
rect 17727 24633 17739 24667
rect 17681 24627 17739 24633
rect 15102 24596 15108 24608
rect 14752 24568 15108 24596
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 17586 24556 17592 24608
rect 17644 24596 17650 24608
rect 17865 24599 17923 24605
rect 17865 24596 17877 24599
rect 17644 24568 17877 24596
rect 17644 24556 17650 24568
rect 17865 24565 17877 24568
rect 17911 24565 17923 24599
rect 17865 24559 17923 24565
rect 1104 24506 18860 24528
rect 1104 24454 3915 24506
rect 3967 24454 3979 24506
rect 4031 24454 4043 24506
rect 4095 24454 4107 24506
rect 4159 24454 4171 24506
rect 4223 24454 9846 24506
rect 9898 24454 9910 24506
rect 9962 24454 9974 24506
rect 10026 24454 10038 24506
rect 10090 24454 10102 24506
rect 10154 24454 15776 24506
rect 15828 24454 15840 24506
rect 15892 24454 15904 24506
rect 15956 24454 15968 24506
rect 16020 24454 16032 24506
rect 16084 24454 18860 24506
rect 1104 24432 18860 24454
rect 5166 24392 5172 24404
rect 5127 24364 5172 24392
rect 5166 24352 5172 24364
rect 5224 24352 5230 24404
rect 14737 24395 14795 24401
rect 14737 24361 14749 24395
rect 14783 24392 14795 24395
rect 15470 24392 15476 24404
rect 14783 24364 15476 24392
rect 14783 24361 14795 24364
rect 14737 24355 14795 24361
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 16577 24395 16635 24401
rect 16577 24361 16589 24395
rect 16623 24392 16635 24395
rect 16758 24392 16764 24404
rect 16623 24364 16764 24392
rect 16623 24361 16635 24364
rect 16577 24355 16635 24361
rect 16758 24352 16764 24364
rect 16816 24352 16822 24404
rect 17126 24392 17132 24404
rect 17087 24364 17132 24392
rect 17126 24352 17132 24364
rect 17184 24352 17190 24404
rect 2406 24216 2412 24268
rect 2464 24256 2470 24268
rect 2501 24259 2559 24265
rect 2501 24256 2513 24259
rect 2464 24228 2513 24256
rect 2464 24216 2470 24228
rect 2501 24225 2513 24228
rect 2547 24256 2559 24259
rect 3789 24259 3847 24265
rect 3789 24256 3801 24259
rect 2547 24228 3801 24256
rect 2547 24225 2559 24228
rect 2501 24219 2559 24225
rect 3789 24225 3801 24228
rect 3835 24256 3847 24259
rect 3878 24256 3884 24268
rect 3835 24228 3884 24256
rect 3835 24225 3847 24228
rect 3789 24219 3847 24225
rect 3878 24216 3884 24228
rect 3936 24216 3942 24268
rect 3973 24259 4031 24265
rect 3973 24225 3985 24259
rect 4019 24256 4031 24259
rect 4338 24256 4344 24268
rect 4019 24228 4344 24256
rect 4019 24225 4031 24228
rect 3973 24219 4031 24225
rect 4338 24216 4344 24228
rect 4396 24256 4402 24268
rect 14369 24259 14427 24265
rect 4396 24228 5304 24256
rect 4396 24216 4402 24228
rect 5276 24197 5304 24228
rect 14369 24225 14381 24259
rect 14415 24256 14427 24259
rect 17862 24256 17868 24268
rect 14415 24228 15332 24256
rect 14415 24225 14427 24228
rect 14369 24219 14427 24225
rect 2593 24191 2651 24197
rect 2593 24157 2605 24191
rect 2639 24157 2651 24191
rect 2593 24151 2651 24157
rect 4065 24191 4123 24197
rect 4065 24157 4077 24191
rect 4111 24157 4123 24191
rect 4065 24151 4123 24157
rect 5261 24191 5319 24197
rect 5261 24157 5273 24191
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 2608 24120 2636 24151
rect 3694 24120 3700 24132
rect 2608 24092 3700 24120
rect 3694 24080 3700 24092
rect 3752 24120 3758 24132
rect 4080 24120 4108 24151
rect 14090 24148 14096 24200
rect 14148 24188 14154 24200
rect 14458 24188 14464 24200
rect 14148 24160 14464 24188
rect 14148 24148 14154 24160
rect 14458 24148 14464 24160
rect 14516 24188 14522 24200
rect 14553 24191 14611 24197
rect 14553 24188 14565 24191
rect 14516 24160 14565 24188
rect 14516 24148 14522 24160
rect 14553 24157 14565 24160
rect 14599 24157 14611 24191
rect 15194 24188 15200 24200
rect 15155 24160 15200 24188
rect 14553 24151 14611 24157
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 15304 24188 15332 24228
rect 16316 24228 17868 24256
rect 16316 24188 16344 24228
rect 17862 24216 17868 24228
rect 17920 24216 17926 24268
rect 15304 24160 16344 24188
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24188 17371 24191
rect 18138 24188 18144 24200
rect 17359 24160 18144 24188
rect 17359 24157 17371 24160
rect 17313 24151 17371 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 3752 24092 4108 24120
rect 12437 24123 12495 24129
rect 3752 24080 3758 24092
rect 12437 24089 12449 24123
rect 12483 24120 12495 24123
rect 15464 24123 15522 24129
rect 12483 24092 15424 24120
rect 12483 24089 12495 24092
rect 12437 24083 12495 24089
rect 2958 24052 2964 24064
rect 2919 24024 2964 24052
rect 2958 24012 2964 24024
rect 3016 24012 3022 24064
rect 3142 24012 3148 24064
rect 3200 24052 3206 24064
rect 3789 24055 3847 24061
rect 3789 24052 3801 24055
rect 3200 24024 3801 24052
rect 3200 24012 3206 24024
rect 3789 24021 3801 24024
rect 3835 24021 3847 24055
rect 3789 24015 3847 24021
rect 10502 24012 10508 24064
rect 10560 24052 10566 24064
rect 11149 24055 11207 24061
rect 11149 24052 11161 24055
rect 10560 24024 11161 24052
rect 10560 24012 10566 24024
rect 11149 24021 11161 24024
rect 11195 24052 11207 24055
rect 11974 24052 11980 24064
rect 11195 24024 11980 24052
rect 11195 24021 11207 24024
rect 11149 24015 11207 24021
rect 11974 24012 11980 24024
rect 12032 24012 12038 24064
rect 15396 24052 15424 24092
rect 15464 24089 15476 24123
rect 15510 24120 15522 24123
rect 15562 24120 15568 24132
rect 15510 24092 15568 24120
rect 15510 24089 15522 24092
rect 15464 24083 15522 24089
rect 15562 24080 15568 24092
rect 15620 24080 15626 24132
rect 16574 24080 16580 24132
rect 16632 24120 16638 24132
rect 17497 24123 17555 24129
rect 17497 24120 17509 24123
rect 16632 24092 17509 24120
rect 16632 24080 16638 24092
rect 17497 24089 17509 24092
rect 17543 24120 17555 24123
rect 17586 24120 17592 24132
rect 17543 24092 17592 24120
rect 17543 24089 17555 24092
rect 17497 24083 17555 24089
rect 17586 24080 17592 24092
rect 17644 24080 17650 24132
rect 17681 24123 17739 24129
rect 17681 24089 17693 24123
rect 17727 24120 17739 24123
rect 18046 24120 18052 24132
rect 17727 24092 18052 24120
rect 17727 24089 17739 24092
rect 17681 24083 17739 24089
rect 18046 24080 18052 24092
rect 18104 24080 18110 24132
rect 16114 24052 16120 24064
rect 15396 24024 16120 24052
rect 16114 24012 16120 24024
rect 16172 24012 16178 24064
rect 17402 24012 17408 24064
rect 17460 24052 17466 24064
rect 17460 24024 17505 24052
rect 17460 24012 17466 24024
rect 1104 23962 18860 23984
rect 1104 23910 6880 23962
rect 6932 23910 6944 23962
rect 6996 23910 7008 23962
rect 7060 23910 7072 23962
rect 7124 23910 7136 23962
rect 7188 23910 12811 23962
rect 12863 23910 12875 23962
rect 12927 23910 12939 23962
rect 12991 23910 13003 23962
rect 13055 23910 13067 23962
rect 13119 23910 18860 23962
rect 1104 23888 18860 23910
rect 3237 23851 3295 23857
rect 3237 23817 3249 23851
rect 3283 23848 3295 23851
rect 4246 23848 4252 23860
rect 3283 23820 4252 23848
rect 3283 23817 3295 23820
rect 3237 23811 3295 23817
rect 4246 23808 4252 23820
rect 4304 23808 4310 23860
rect 17402 23808 17408 23860
rect 17460 23848 17466 23860
rect 18141 23851 18199 23857
rect 18141 23848 18153 23851
rect 17460 23820 18153 23848
rect 17460 23808 17466 23820
rect 18141 23817 18153 23820
rect 18187 23817 18199 23851
rect 18141 23811 18199 23817
rect 3878 23780 3884 23792
rect 3839 23752 3884 23780
rect 3878 23740 3884 23752
rect 3936 23740 3942 23792
rect 12250 23740 12256 23792
rect 12308 23780 12314 23792
rect 15194 23780 15200 23792
rect 12308 23752 15200 23780
rect 12308 23740 12314 23752
rect 2958 23712 2964 23724
rect 2919 23684 2964 23712
rect 2958 23672 2964 23684
rect 3016 23672 3022 23724
rect 3145 23715 3203 23721
rect 3145 23681 3157 23715
rect 3191 23712 3203 23715
rect 3234 23712 3240 23724
rect 3191 23684 3240 23712
rect 3191 23681 3203 23684
rect 3145 23675 3203 23681
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 3694 23672 3700 23724
rect 3752 23712 3758 23724
rect 4065 23715 4123 23721
rect 4065 23712 4077 23715
rect 3752 23684 4077 23712
rect 3752 23672 3758 23684
rect 4065 23681 4077 23684
rect 4111 23681 4123 23715
rect 7190 23712 7196 23724
rect 7151 23684 7196 23712
rect 4065 23675 4123 23681
rect 7190 23672 7196 23684
rect 7248 23672 7254 23724
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 7300 23684 7665 23712
rect 7300 23656 7328 23684
rect 7653 23681 7665 23684
rect 7699 23681 7711 23715
rect 7653 23675 7711 23681
rect 7837 23715 7895 23721
rect 7837 23681 7849 23715
rect 7883 23712 7895 23715
rect 8202 23712 8208 23724
rect 7883 23684 8208 23712
rect 7883 23681 7895 23684
rect 7837 23675 7895 23681
rect 8202 23672 8208 23684
rect 8260 23672 8266 23724
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13311 23684 13768 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 6730 23604 6736 23656
rect 6788 23644 6794 23656
rect 7282 23644 7288 23656
rect 6788 23616 7288 23644
rect 6788 23604 6794 23616
rect 7282 23604 7288 23616
rect 7340 23604 7346 23656
rect 13096 23644 13124 23675
rect 13630 23644 13636 23656
rect 13096 23616 13636 23644
rect 13630 23604 13636 23616
rect 13688 23604 13694 23656
rect 8110 23576 8116 23588
rect 7576 23548 8116 23576
rect 7576 23520 7604 23548
rect 8110 23536 8116 23548
rect 8168 23536 8174 23588
rect 3418 23508 3424 23520
rect 3379 23480 3424 23508
rect 3418 23468 3424 23480
rect 3476 23468 3482 23520
rect 7009 23511 7067 23517
rect 7009 23477 7021 23511
rect 7055 23508 7067 23511
rect 7558 23508 7564 23520
rect 7055 23480 7564 23508
rect 7055 23477 7067 23480
rect 7009 23471 7067 23477
rect 7558 23468 7564 23480
rect 7616 23468 7622 23520
rect 7834 23508 7840 23520
rect 7795 23480 7840 23508
rect 7834 23468 7840 23480
rect 7892 23468 7898 23520
rect 13262 23508 13268 23520
rect 13223 23480 13268 23508
rect 13262 23468 13268 23480
rect 13320 23468 13326 23520
rect 13740 23517 13768 23684
rect 14826 23672 14832 23724
rect 14884 23721 14890 23724
rect 15120 23721 15148 23752
rect 15194 23740 15200 23752
rect 15252 23780 15258 23792
rect 15252 23752 16804 23780
rect 15252 23740 15258 23752
rect 16776 23724 16804 23752
rect 14884 23712 14896 23721
rect 15105 23715 15163 23721
rect 14884 23684 14929 23712
rect 14884 23675 14896 23684
rect 15105 23681 15117 23715
rect 15151 23681 15163 23715
rect 16114 23712 16120 23724
rect 16075 23684 16120 23712
rect 15105 23675 15163 23681
rect 14884 23672 14890 23675
rect 16114 23672 16120 23684
rect 16172 23672 16178 23724
rect 16758 23712 16764 23724
rect 16671 23684 16764 23712
rect 16758 23672 16764 23684
rect 16816 23672 16822 23724
rect 17028 23715 17086 23721
rect 17028 23681 17040 23715
rect 17074 23712 17086 23715
rect 17586 23712 17592 23724
rect 17074 23684 17592 23712
rect 17074 23681 17086 23684
rect 17028 23675 17086 23681
rect 17586 23672 17592 23684
rect 17644 23672 17650 23724
rect 13725 23511 13783 23517
rect 13725 23477 13737 23511
rect 13771 23508 13783 23511
rect 13814 23508 13820 23520
rect 13771 23480 13820 23508
rect 13771 23477 13783 23480
rect 13725 23471 13783 23477
rect 13814 23468 13820 23480
rect 13872 23468 13878 23520
rect 15933 23511 15991 23517
rect 15933 23477 15945 23511
rect 15979 23508 15991 23511
rect 16206 23508 16212 23520
rect 15979 23480 16212 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 1104 23418 18860 23440
rect 1104 23366 3915 23418
rect 3967 23366 3979 23418
rect 4031 23366 4043 23418
rect 4095 23366 4107 23418
rect 4159 23366 4171 23418
rect 4223 23366 9846 23418
rect 9898 23366 9910 23418
rect 9962 23366 9974 23418
rect 10026 23366 10038 23418
rect 10090 23366 10102 23418
rect 10154 23366 15776 23418
rect 15828 23366 15840 23418
rect 15892 23366 15904 23418
rect 15956 23366 15968 23418
rect 16020 23366 16032 23418
rect 16084 23366 18860 23418
rect 1104 23344 18860 23366
rect 2685 23307 2743 23313
rect 2685 23273 2697 23307
rect 2731 23304 2743 23307
rect 3326 23304 3332 23316
rect 2731 23276 3332 23304
rect 2731 23273 2743 23276
rect 2685 23267 2743 23273
rect 3326 23264 3332 23276
rect 3384 23264 3390 23316
rect 3418 23264 3424 23316
rect 3476 23304 3482 23316
rect 3789 23307 3847 23313
rect 3789 23304 3801 23307
rect 3476 23276 3801 23304
rect 3476 23264 3482 23276
rect 3789 23273 3801 23276
rect 3835 23273 3847 23307
rect 3789 23267 3847 23273
rect 5537 23307 5595 23313
rect 5537 23273 5549 23307
rect 5583 23304 5595 23307
rect 5718 23304 5724 23316
rect 5583 23276 5724 23304
rect 5583 23273 5595 23276
rect 5537 23267 5595 23273
rect 5718 23264 5724 23276
rect 5776 23304 5782 23316
rect 9122 23304 9128 23316
rect 5776 23276 6224 23304
rect 9083 23276 9128 23304
rect 5776 23264 5782 23276
rect 2958 23196 2964 23248
rect 3016 23236 3022 23248
rect 3053 23239 3111 23245
rect 3053 23236 3065 23239
rect 3016 23208 3065 23236
rect 3016 23196 3022 23208
rect 3053 23205 3065 23208
rect 3099 23236 3111 23239
rect 6089 23239 6147 23245
rect 3099 23208 4108 23236
rect 3099 23205 3111 23208
rect 3053 23199 3111 23205
rect 3234 23128 3240 23180
rect 3292 23168 3298 23180
rect 4080 23177 4108 23208
rect 6089 23205 6101 23239
rect 6135 23205 6147 23239
rect 6089 23199 6147 23205
rect 3973 23171 4031 23177
rect 3973 23168 3985 23171
rect 3292 23140 3985 23168
rect 3292 23128 3298 23140
rect 3973 23137 3985 23140
rect 4019 23137 4031 23171
rect 3973 23131 4031 23137
rect 4065 23171 4123 23177
rect 4065 23137 4077 23171
rect 4111 23137 4123 23171
rect 6104 23168 6132 23199
rect 4065 23131 4123 23137
rect 5368 23140 6132 23168
rect 2866 23100 2872 23112
rect 2827 23072 2872 23100
rect 2866 23060 2872 23072
rect 2924 23060 2930 23112
rect 2958 23060 2964 23112
rect 3016 23100 3022 23112
rect 3016 23072 3061 23100
rect 3016 23060 3022 23072
rect 3142 23060 3148 23112
rect 3200 23100 3206 23112
rect 5368 23109 5396 23140
rect 5353 23103 5411 23109
rect 3200 23072 3245 23100
rect 3200 23060 3206 23072
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 5626 23060 5632 23112
rect 5684 23100 5690 23112
rect 6196 23100 6224 23276
rect 9122 23264 9128 23276
rect 9180 23264 9186 23316
rect 8941 23239 8999 23245
rect 8941 23205 8953 23239
rect 8987 23205 8999 23239
rect 8941 23199 8999 23205
rect 6365 23103 6423 23109
rect 6365 23100 6377 23103
rect 5684 23072 6040 23100
rect 6196 23072 6377 23100
rect 5684 23060 5690 23072
rect 6012 22976 6040 23072
rect 6365 23069 6377 23072
rect 6411 23100 6423 23103
rect 6454 23100 6460 23112
rect 6411 23072 6460 23100
rect 6411 23069 6423 23072
rect 6365 23063 6423 23069
rect 6454 23060 6460 23072
rect 6512 23060 6518 23112
rect 7009 23103 7067 23109
rect 7009 23069 7021 23103
rect 7055 23100 7067 23103
rect 7282 23100 7288 23112
rect 7055 23072 7288 23100
rect 7055 23069 7067 23072
rect 7009 23063 7067 23069
rect 7282 23060 7288 23072
rect 7340 23060 7346 23112
rect 8294 23100 8300 23112
rect 8255 23072 8300 23100
rect 8294 23060 8300 23072
rect 8352 23060 8358 23112
rect 8389 23103 8447 23109
rect 8389 23069 8401 23103
rect 8435 23100 8447 23103
rect 8956 23100 8984 23199
rect 13630 23196 13636 23248
rect 13688 23236 13694 23248
rect 14277 23239 14335 23245
rect 13688 23208 14228 23236
rect 13688 23196 13694 23208
rect 13446 23168 13452 23180
rect 13407 23140 13452 23168
rect 13446 23128 13452 23140
rect 13504 23168 13510 23180
rect 14093 23171 14151 23177
rect 14093 23168 14105 23171
rect 13504 23140 14105 23168
rect 13504 23128 13510 23140
rect 14093 23137 14105 23140
rect 14139 23137 14151 23171
rect 14200 23168 14228 23208
rect 14277 23205 14289 23239
rect 14323 23236 14335 23239
rect 14550 23236 14556 23248
rect 14323 23208 14556 23236
rect 14323 23205 14335 23208
rect 14277 23199 14335 23205
rect 14550 23196 14556 23208
rect 14608 23196 14614 23248
rect 15381 23171 15439 23177
rect 15381 23168 15393 23171
rect 14200 23140 15393 23168
rect 14093 23131 14151 23137
rect 15381 23137 15393 23140
rect 15427 23137 15439 23171
rect 15381 23131 15439 23137
rect 15933 23171 15991 23177
rect 15933 23137 15945 23171
rect 15979 23168 15991 23171
rect 16574 23168 16580 23180
rect 15979 23140 16580 23168
rect 15979 23137 15991 23140
rect 15933 23131 15991 23137
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 16758 23168 16764 23180
rect 16719 23140 16764 23168
rect 16758 23128 16764 23140
rect 16816 23128 16822 23180
rect 10226 23100 10232 23112
rect 8435 23072 10232 23100
rect 8435 23069 8447 23072
rect 8389 23063 8447 23069
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 13170 23100 13176 23112
rect 13131 23072 13176 23100
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 13262 23060 13268 23112
rect 13320 23100 13326 23112
rect 13541 23103 13599 23109
rect 13320 23072 13365 23100
rect 13320 23060 13326 23072
rect 13541 23069 13553 23103
rect 13587 23069 13599 23103
rect 13541 23063 13599 23069
rect 6086 22992 6092 23044
rect 6144 23032 6150 23044
rect 7377 23035 7435 23041
rect 6144 23004 6189 23032
rect 6144 22992 6150 23004
rect 7377 23001 7389 23035
rect 7423 23032 7435 23035
rect 8113 23035 8171 23041
rect 8113 23032 8125 23035
rect 7423 23004 8125 23032
rect 7423 23001 7435 23004
rect 7377 22995 7435 23001
rect 8113 23001 8125 23004
rect 8159 23001 8171 23035
rect 8113 22995 8171 23001
rect 4433 22967 4491 22973
rect 4433 22933 4445 22967
rect 4479 22964 4491 22967
rect 4706 22964 4712 22976
rect 4479 22936 4712 22964
rect 4479 22933 4491 22936
rect 4433 22927 4491 22933
rect 4706 22924 4712 22936
rect 4764 22924 4770 22976
rect 5166 22964 5172 22976
rect 5127 22936 5172 22964
rect 5166 22924 5172 22936
rect 5224 22924 5230 22976
rect 5994 22924 6000 22976
rect 6052 22964 6058 22976
rect 6273 22967 6331 22973
rect 6273 22964 6285 22967
rect 6052 22936 6285 22964
rect 6052 22924 6058 22936
rect 6273 22933 6285 22936
rect 6319 22933 6331 22967
rect 6273 22927 6331 22933
rect 6362 22924 6368 22976
rect 6420 22964 6426 22976
rect 7392 22964 7420 22995
rect 8202 22992 8208 23044
rect 8260 23032 8266 23044
rect 9093 23035 9151 23041
rect 9093 23032 9105 23035
rect 8260 23004 9105 23032
rect 8260 22992 8266 23004
rect 9093 23001 9105 23004
rect 9139 23032 9151 23035
rect 9306 23032 9312 23044
rect 9139 23001 9168 23032
rect 9267 23004 9312 23032
rect 9093 22995 9168 23001
rect 8386 22964 8392 22976
rect 6420 22936 7420 22964
rect 8347 22936 8392 22964
rect 6420 22924 6426 22936
rect 8386 22924 8392 22936
rect 8444 22924 8450 22976
rect 9140 22964 9168 22995
rect 9306 22992 9312 23004
rect 9364 22992 9370 23044
rect 13556 22976 13584 23063
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 15197 23103 15255 23109
rect 15197 23100 15209 23103
rect 13872 23072 15209 23100
rect 13872 23060 13878 23072
rect 15197 23069 15209 23072
rect 15243 23069 15255 23103
rect 15197 23063 15255 23069
rect 16022 23060 16028 23112
rect 16080 23100 16086 23112
rect 16117 23103 16175 23109
rect 16117 23100 16129 23103
rect 16080 23072 16129 23100
rect 16080 23060 16086 23072
rect 16117 23069 16129 23072
rect 16163 23069 16175 23103
rect 16117 23063 16175 23069
rect 14553 23035 14611 23041
rect 14553 23001 14565 23035
rect 14599 23032 14611 23035
rect 14642 23032 14648 23044
rect 14599 23004 14648 23032
rect 14599 23001 14611 23004
rect 14553 22995 14611 23001
rect 14642 22992 14648 23004
rect 14700 22992 14706 23044
rect 17028 23035 17086 23041
rect 17028 23001 17040 23035
rect 17074 23032 17086 23035
rect 17126 23032 17132 23044
rect 17074 23004 17132 23032
rect 17074 23001 17086 23004
rect 17028 22995 17086 23001
rect 17126 22992 17132 23004
rect 17184 22992 17190 23044
rect 10502 22964 10508 22976
rect 9140 22936 10508 22964
rect 10502 22924 10508 22936
rect 10560 22924 10566 22976
rect 12618 22924 12624 22976
rect 12676 22964 12682 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12676 22936 13001 22964
rect 12676 22924 12682 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 13538 22964 13544 22976
rect 13451 22936 13544 22964
rect 12989 22927 13047 22933
rect 13538 22924 13544 22936
rect 13596 22964 13602 22976
rect 15013 22967 15071 22973
rect 15013 22964 15025 22967
rect 13596 22936 15025 22964
rect 13596 22924 13602 22936
rect 15013 22933 15025 22936
rect 15059 22933 15071 22967
rect 15013 22927 15071 22933
rect 16301 22967 16359 22973
rect 16301 22933 16313 22967
rect 16347 22964 16359 22967
rect 16942 22964 16948 22976
rect 16347 22936 16948 22964
rect 16347 22933 16359 22936
rect 16301 22927 16359 22933
rect 16942 22924 16948 22936
rect 17000 22924 17006 22976
rect 18046 22924 18052 22976
rect 18104 22964 18110 22976
rect 18141 22967 18199 22973
rect 18141 22964 18153 22967
rect 18104 22936 18153 22964
rect 18104 22924 18110 22936
rect 18141 22933 18153 22936
rect 18187 22933 18199 22967
rect 18141 22927 18199 22933
rect 1104 22874 18860 22896
rect 1104 22822 6880 22874
rect 6932 22822 6944 22874
rect 6996 22822 7008 22874
rect 7060 22822 7072 22874
rect 7124 22822 7136 22874
rect 7188 22822 12811 22874
rect 12863 22822 12875 22874
rect 12927 22822 12939 22874
rect 12991 22822 13003 22874
rect 13055 22822 13067 22874
rect 13119 22822 18860 22874
rect 1104 22800 18860 22822
rect 3234 22760 3240 22772
rect 3195 22732 3240 22760
rect 3234 22720 3240 22732
rect 3292 22720 3298 22772
rect 3786 22760 3792 22772
rect 3747 22732 3792 22760
rect 3786 22720 3792 22732
rect 3844 22720 3850 22772
rect 4706 22760 4712 22772
rect 3896 22732 4712 22760
rect 3896 22701 3924 22732
rect 4706 22720 4712 22732
rect 4764 22720 4770 22772
rect 5442 22720 5448 22772
rect 5500 22760 5506 22772
rect 6362 22760 6368 22772
rect 5500 22732 6368 22760
rect 5500 22720 5506 22732
rect 6362 22720 6368 22732
rect 6420 22720 6426 22772
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 10327 22763 10385 22769
rect 10327 22760 10339 22763
rect 8352 22732 10339 22760
rect 8352 22720 8358 22732
rect 10327 22729 10339 22732
rect 10373 22729 10385 22763
rect 10327 22723 10385 22729
rect 13170 22720 13176 22772
rect 13228 22760 13234 22772
rect 14093 22763 14151 22769
rect 14093 22760 14105 22763
rect 13228 22732 14105 22760
rect 13228 22720 13234 22732
rect 14093 22729 14105 22732
rect 14139 22729 14151 22763
rect 14093 22723 14151 22729
rect 3881 22695 3939 22701
rect 3881 22661 3893 22695
rect 3927 22661 3939 22695
rect 3881 22655 3939 22661
rect 4448 22664 8340 22692
rect 4448 22636 4476 22664
rect 2866 22584 2872 22636
rect 2924 22624 2930 22636
rect 2961 22627 3019 22633
rect 2961 22624 2973 22627
rect 2924 22596 2973 22624
rect 2924 22584 2930 22596
rect 2961 22593 2973 22596
rect 3007 22624 3019 22627
rect 3326 22624 3332 22636
rect 3007 22596 3332 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 3326 22584 3332 22596
rect 3384 22584 3390 22636
rect 4430 22624 4436 22636
rect 4343 22596 4436 22624
rect 4430 22584 4436 22596
rect 4488 22584 4494 22636
rect 4700 22627 4758 22633
rect 4700 22593 4712 22627
rect 4746 22624 4758 22627
rect 5166 22624 5172 22636
rect 4746 22596 5172 22624
rect 4746 22593 4758 22596
rect 4700 22587 4758 22593
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7650 22624 7656 22636
rect 6963 22596 7656 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 8312 22568 8340 22664
rect 8386 22652 8392 22704
rect 8444 22692 8450 22704
rect 8634 22695 8692 22701
rect 8634 22692 8646 22695
rect 8444 22664 8646 22692
rect 8444 22652 8450 22664
rect 8634 22661 8646 22664
rect 8680 22661 8692 22695
rect 8634 22655 8692 22661
rect 9122 22652 9128 22704
rect 9180 22692 9186 22704
rect 10413 22695 10471 22701
rect 10413 22692 10425 22695
rect 9180 22664 10425 22692
rect 9180 22652 9186 22664
rect 10413 22661 10425 22664
rect 10459 22661 10471 22695
rect 10413 22655 10471 22661
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 9784 22596 10241 22624
rect 3234 22556 3240 22568
rect 3195 22528 3240 22556
rect 3234 22516 3240 22528
rect 3292 22516 3298 22568
rect 7193 22559 7251 22565
rect 7193 22525 7205 22559
rect 7239 22556 7251 22559
rect 7374 22556 7380 22568
rect 7239 22528 7380 22556
rect 7239 22525 7251 22528
rect 7193 22519 7251 22525
rect 7374 22516 7380 22528
rect 7432 22516 7438 22568
rect 8294 22516 8300 22568
rect 8352 22556 8358 22568
rect 8389 22559 8447 22565
rect 8389 22556 8401 22559
rect 8352 22528 8401 22556
rect 8352 22516 8358 22528
rect 8389 22525 8401 22528
rect 8435 22525 8447 22559
rect 8389 22519 8447 22525
rect 2958 22448 2964 22500
rect 3016 22488 3022 22500
rect 3053 22491 3111 22497
rect 3053 22488 3065 22491
rect 3016 22460 3065 22488
rect 3016 22448 3022 22460
rect 3053 22457 3065 22460
rect 3099 22457 3111 22491
rect 3053 22451 3111 22457
rect 5718 22380 5724 22432
rect 5776 22420 5782 22432
rect 5813 22423 5871 22429
rect 5813 22420 5825 22423
rect 5776 22392 5825 22420
rect 5776 22380 5782 22392
rect 5813 22389 5825 22392
rect 5859 22389 5871 22423
rect 5813 22383 5871 22389
rect 9030 22380 9036 22432
rect 9088 22420 9094 22432
rect 9306 22420 9312 22432
rect 9088 22392 9312 22420
rect 9088 22380 9094 22392
rect 9306 22380 9312 22392
rect 9364 22420 9370 22432
rect 9784 22429 9812 22596
rect 10229 22593 10241 22596
rect 10275 22593 10287 22627
rect 10502 22624 10508 22636
rect 10463 22596 10508 22624
rect 10229 22587 10287 22593
rect 10502 22584 10508 22596
rect 10560 22584 10566 22636
rect 11514 22624 11520 22636
rect 11475 22596 11520 22624
rect 11514 22584 11520 22596
rect 11572 22584 11578 22636
rect 12526 22633 12532 22636
rect 12520 22587 12532 22633
rect 12584 22624 12590 22636
rect 15010 22624 15016 22636
rect 12584 22596 12620 22624
rect 14971 22596 15016 22624
rect 12526 22584 12532 22587
rect 12584 22584 12590 22596
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22624 15347 22627
rect 15654 22624 15660 22636
rect 15335 22596 15660 22624
rect 15335 22593 15347 22596
rect 15289 22587 15347 22593
rect 15654 22584 15660 22596
rect 15712 22624 15718 22636
rect 16022 22624 16028 22636
rect 15712 22596 16028 22624
rect 15712 22584 15718 22596
rect 16022 22584 16028 22596
rect 16080 22584 16086 22636
rect 16669 22627 16727 22633
rect 16669 22593 16681 22627
rect 16715 22624 16727 22627
rect 16758 22624 16764 22636
rect 16715 22596 16764 22624
rect 16715 22593 16727 22596
rect 16669 22587 16727 22593
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 16942 22633 16948 22636
rect 16936 22587 16948 22633
rect 17000 22624 17006 22636
rect 17000 22596 17036 22624
rect 16942 22584 16948 22587
rect 17000 22584 17006 22596
rect 11238 22516 11244 22568
rect 11296 22556 11302 22568
rect 12250 22556 12256 22568
rect 11296 22528 12256 22556
rect 11296 22516 11302 22528
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 14550 22556 14556 22568
rect 14511 22528 14556 22556
rect 14550 22516 14556 22528
rect 14608 22516 14614 22568
rect 13630 22488 13636 22500
rect 13591 22460 13636 22488
rect 13630 22448 13636 22460
rect 13688 22448 13694 22500
rect 14277 22491 14335 22497
rect 14277 22457 14289 22491
rect 14323 22488 14335 22491
rect 14642 22488 14648 22500
rect 14323 22460 14648 22488
rect 14323 22457 14335 22460
rect 14277 22451 14335 22457
rect 14642 22448 14648 22460
rect 14700 22448 14706 22500
rect 9769 22423 9827 22429
rect 9769 22420 9781 22423
rect 9364 22392 9781 22420
rect 9364 22380 9370 22392
rect 9769 22389 9781 22392
rect 9815 22389 9827 22423
rect 9769 22383 9827 22389
rect 11606 22380 11612 22432
rect 11664 22420 11670 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 11664 22392 11713 22420
rect 11664 22380 11670 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 18049 22423 18107 22429
rect 18049 22389 18061 22423
rect 18095 22420 18107 22423
rect 18138 22420 18144 22432
rect 18095 22392 18144 22420
rect 18095 22389 18107 22392
rect 18049 22383 18107 22389
rect 18138 22380 18144 22392
rect 18196 22380 18202 22432
rect 1104 22330 18860 22352
rect 1104 22278 3915 22330
rect 3967 22278 3979 22330
rect 4031 22278 4043 22330
rect 4095 22278 4107 22330
rect 4159 22278 4171 22330
rect 4223 22278 9846 22330
rect 9898 22278 9910 22330
rect 9962 22278 9974 22330
rect 10026 22278 10038 22330
rect 10090 22278 10102 22330
rect 10154 22278 15776 22330
rect 15828 22278 15840 22330
rect 15892 22278 15904 22330
rect 15956 22278 15968 22330
rect 16020 22278 16032 22330
rect 16084 22278 18860 22330
rect 1104 22256 18860 22278
rect 2774 22176 2780 22228
rect 2832 22216 2838 22228
rect 3145 22219 3203 22225
rect 3145 22216 3157 22219
rect 2832 22188 3157 22216
rect 2832 22176 2838 22188
rect 3145 22185 3157 22188
rect 3191 22216 3203 22219
rect 3234 22216 3240 22228
rect 3191 22188 3240 22216
rect 3191 22185 3203 22188
rect 3145 22179 3203 22185
rect 3234 22176 3240 22188
rect 3292 22176 3298 22228
rect 7650 22176 7656 22228
rect 7708 22216 7714 22228
rect 7708 22188 12434 22216
rect 7708 22176 7714 22188
rect 12406 22148 12434 22188
rect 13262 22176 13268 22228
rect 13320 22216 13326 22228
rect 13449 22219 13507 22225
rect 13449 22216 13461 22219
rect 13320 22188 13461 22216
rect 13320 22176 13326 22188
rect 13449 22185 13461 22188
rect 13495 22185 13507 22219
rect 13449 22179 13507 22185
rect 13354 22148 13360 22160
rect 12406 22120 13360 22148
rect 13354 22108 13360 22120
rect 13412 22108 13418 22160
rect 3881 22083 3939 22089
rect 3881 22080 3893 22083
rect 2424 22052 3893 22080
rect 2424 22021 2452 22052
rect 3881 22049 3893 22052
rect 3927 22049 3939 22083
rect 5718 22080 5724 22092
rect 5679 22052 5724 22080
rect 3881 22043 3939 22049
rect 5718 22040 5724 22052
rect 5776 22040 5782 22092
rect 5994 22080 6000 22092
rect 5955 22052 6000 22080
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 9585 22083 9643 22089
rect 9585 22080 9597 22083
rect 8312 22052 9597 22080
rect 8312 22024 8340 22052
rect 9585 22049 9597 22052
rect 9631 22049 9643 22083
rect 9585 22043 9643 22049
rect 10686 22040 10692 22092
rect 10744 22080 10750 22092
rect 13446 22080 13452 22092
rect 10744 22052 11652 22080
rect 10744 22040 10750 22052
rect 2409 22015 2467 22021
rect 2409 21981 2421 22015
rect 2455 21981 2467 22015
rect 2409 21975 2467 21981
rect 2593 22015 2651 22021
rect 2593 21981 2605 22015
rect 2639 22012 2651 22015
rect 2774 22012 2780 22024
rect 2639 21984 2780 22012
rect 2639 21981 2651 21984
rect 2593 21975 2651 21981
rect 2774 21972 2780 21984
rect 2832 21972 2838 22024
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 21981 3111 22015
rect 3053 21975 3111 21981
rect 3237 22015 3295 22021
rect 3237 21981 3249 22015
rect 3283 22012 3295 22015
rect 3694 22012 3700 22024
rect 3283 21984 3700 22012
rect 3283 21981 3295 21984
rect 3237 21975 3295 21981
rect 3068 21944 3096 21975
rect 3694 21972 3700 21984
rect 3752 21972 3758 22024
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 22012 4123 22015
rect 4338 22012 4344 22024
rect 4111 21984 4344 22012
rect 4111 21981 4123 21984
rect 4065 21975 4123 21981
rect 4080 21944 4108 21975
rect 4338 21972 4344 21984
rect 4396 22012 4402 22024
rect 4522 22012 4528 22024
rect 4396 21984 4528 22012
rect 4396 21972 4402 21984
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 5261 22015 5319 22021
rect 5261 21981 5273 22015
rect 5307 21981 5319 22015
rect 5261 21975 5319 21981
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 22012 7067 22015
rect 8294 22012 8300 22024
rect 7055 21984 8300 22012
rect 7055 21981 7067 21984
rect 7009 21975 7067 21981
rect 3068 21916 4108 21944
rect 4249 21947 4307 21953
rect 4249 21913 4261 21947
rect 4295 21913 4307 21947
rect 5276 21944 5304 21975
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 9122 22012 9128 22024
rect 9035 21984 9128 22012
rect 9122 21972 9128 21984
rect 9180 22012 9186 22024
rect 11422 22012 11428 22024
rect 9180 21984 9628 22012
rect 11383 21984 11428 22012
rect 9180 21972 9186 21984
rect 9600 21956 9628 21984
rect 11422 21972 11428 21984
rect 11480 21972 11486 22024
rect 11624 22021 11652 22052
rect 13188 22052 13452 22080
rect 13188 22021 13216 22052
rect 13446 22040 13452 22052
rect 13504 22040 13510 22092
rect 13538 22040 13544 22092
rect 13596 22080 13602 22092
rect 15654 22080 15660 22092
rect 13596 22052 13641 22080
rect 14476 22052 15660 22080
rect 13596 22040 13602 22052
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 13173 22015 13231 22021
rect 13173 21981 13185 22015
rect 13219 21981 13231 22015
rect 13173 21975 13231 21981
rect 13262 21972 13268 22024
rect 13320 22012 13326 22024
rect 14476 22021 14504 22052
rect 15654 22040 15660 22052
rect 15712 22080 15718 22092
rect 17957 22083 18015 22089
rect 15712 22052 17816 22080
rect 15712 22040 15718 22052
rect 14461 22015 14519 22021
rect 13320 21984 13365 22012
rect 13320 21972 13326 21984
rect 14461 21981 14473 22015
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 14550 21972 14556 22024
rect 14608 22012 14614 22024
rect 16960 22021 16988 22052
rect 17788 22021 17816 22052
rect 17957 22049 17969 22083
rect 18003 22080 18015 22083
rect 18138 22080 18144 22092
rect 18003 22052 18144 22080
rect 18003 22049 18015 22052
rect 17957 22043 18015 22049
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 16117 22015 16175 22021
rect 14608 21984 14653 22012
rect 14608 21972 14614 21984
rect 16117 21981 16129 22015
rect 16163 22012 16175 22015
rect 16761 22015 16819 22021
rect 16761 22012 16773 22015
rect 16163 21984 16773 22012
rect 16163 21981 16175 21984
rect 16117 21975 16175 21981
rect 16761 21981 16773 21984
rect 16807 21981 16819 22015
rect 16761 21975 16819 21981
rect 16945 22015 17003 22021
rect 16945 21981 16957 22015
rect 16991 21981 17003 22015
rect 16945 21975 17003 21981
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 21981 17187 22015
rect 17129 21975 17187 21981
rect 17773 22015 17831 22021
rect 17773 21981 17785 22015
rect 17819 21981 17831 22015
rect 17773 21975 17831 21981
rect 7276 21947 7334 21953
rect 5276 21916 7236 21944
rect 4249 21907 4307 21913
rect 2593 21879 2651 21885
rect 2593 21845 2605 21879
rect 2639 21876 2651 21879
rect 2774 21876 2780 21888
rect 2639 21848 2780 21876
rect 2639 21845 2651 21848
rect 2593 21839 2651 21845
rect 2774 21836 2780 21848
rect 2832 21876 2838 21888
rect 2958 21876 2964 21888
rect 2832 21848 2964 21876
rect 2832 21836 2838 21848
rect 2958 21836 2964 21848
rect 3016 21836 3022 21888
rect 3694 21836 3700 21888
rect 3752 21876 3758 21888
rect 4264 21876 4292 21907
rect 4338 21876 4344 21888
rect 3752 21848 4344 21876
rect 3752 21836 3758 21848
rect 4338 21836 4344 21848
rect 4396 21836 4402 21888
rect 5077 21879 5135 21885
rect 5077 21845 5089 21879
rect 5123 21876 5135 21879
rect 5626 21876 5632 21888
rect 5123 21848 5632 21876
rect 5123 21845 5135 21848
rect 5077 21839 5135 21845
rect 5626 21836 5632 21848
rect 5684 21876 5690 21888
rect 6730 21876 6736 21888
rect 5684 21848 6736 21876
rect 5684 21836 5690 21848
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 7208 21876 7236 21916
rect 7276 21913 7288 21947
rect 7322 21944 7334 21947
rect 7834 21944 7840 21956
rect 7322 21916 7840 21944
rect 7322 21913 7334 21916
rect 7276 21907 7334 21913
rect 7834 21904 7840 21916
rect 7892 21904 7898 21956
rect 9582 21904 9588 21956
rect 9640 21904 9646 21956
rect 9852 21947 9910 21953
rect 9852 21913 9864 21947
rect 9898 21944 9910 21947
rect 11517 21947 11575 21953
rect 11517 21944 11529 21947
rect 9898 21916 11529 21944
rect 9898 21913 9910 21916
rect 9852 21907 9910 21913
rect 11517 21913 11529 21916
rect 11563 21913 11575 21947
rect 11517 21907 11575 21913
rect 12989 21947 13047 21953
rect 12989 21913 13001 21947
rect 13035 21944 13047 21947
rect 13538 21944 13544 21956
rect 13035 21916 13544 21944
rect 13035 21913 13047 21916
rect 12989 21907 13047 21913
rect 13538 21904 13544 21916
rect 13596 21904 13602 21956
rect 17144 21944 17172 21975
rect 18046 21944 18052 21956
rect 17144 21916 18052 21944
rect 18046 21904 18052 21916
rect 18104 21904 18110 21956
rect 7374 21876 7380 21888
rect 7208 21848 7380 21876
rect 7374 21836 7380 21848
rect 7432 21836 7438 21888
rect 8110 21836 8116 21888
rect 8168 21876 8174 21888
rect 8389 21879 8447 21885
rect 8389 21876 8401 21879
rect 8168 21848 8401 21876
rect 8168 21836 8174 21848
rect 8389 21845 8401 21848
rect 8435 21845 8447 21879
rect 8389 21839 8447 21845
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 9033 21879 9091 21885
rect 9033 21876 9045 21879
rect 8628 21848 9045 21876
rect 8628 21836 8634 21848
rect 9033 21845 9045 21848
rect 9079 21845 9091 21879
rect 10962 21876 10968 21888
rect 10923 21848 10968 21876
rect 9033 21839 9091 21845
rect 10962 21836 10968 21848
rect 11020 21836 11026 21888
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13504 21848 14289 21876
rect 13504 21836 13510 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 14277 21839 14335 21845
rect 16301 21879 16359 21885
rect 16301 21845 16313 21879
rect 16347 21876 16359 21879
rect 16758 21876 16764 21888
rect 16347 21848 16764 21876
rect 16347 21845 16359 21848
rect 16301 21839 16359 21845
rect 16758 21836 16764 21848
rect 16816 21836 16822 21888
rect 17589 21879 17647 21885
rect 17589 21845 17601 21879
rect 17635 21876 17647 21879
rect 17770 21876 17776 21888
rect 17635 21848 17776 21876
rect 17635 21845 17647 21848
rect 17589 21839 17647 21845
rect 17770 21836 17776 21848
rect 17828 21836 17834 21888
rect 1104 21786 18860 21808
rect 1104 21734 6880 21786
rect 6932 21734 6944 21786
rect 6996 21734 7008 21786
rect 7060 21734 7072 21786
rect 7124 21734 7136 21786
rect 7188 21734 12811 21786
rect 12863 21734 12875 21786
rect 12927 21734 12939 21786
rect 12991 21734 13003 21786
rect 13055 21734 13067 21786
rect 13119 21734 18860 21786
rect 1104 21712 18860 21734
rect 4614 21672 4620 21684
rect 4172 21644 4620 21672
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 2958 21536 2964 21548
rect 2915 21508 2964 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 2958 21496 2964 21508
rect 3016 21536 3022 21548
rect 3326 21536 3332 21548
rect 3016 21508 3332 21536
rect 3016 21496 3022 21508
rect 3326 21496 3332 21508
rect 3384 21496 3390 21548
rect 4172 21545 4200 21644
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 5810 21672 5816 21684
rect 5771 21644 5816 21672
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 10413 21675 10471 21681
rect 10413 21641 10425 21675
rect 10459 21672 10471 21675
rect 10686 21672 10692 21684
rect 10459 21644 10692 21672
rect 10459 21641 10471 21644
rect 10413 21635 10471 21641
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 12526 21632 12532 21684
rect 12584 21672 12590 21684
rect 13265 21675 13323 21681
rect 13265 21672 13277 21675
rect 12584 21644 13277 21672
rect 12584 21632 12590 21644
rect 13265 21641 13277 21644
rect 13311 21641 13323 21675
rect 17126 21672 17132 21684
rect 17087 21644 17132 21672
rect 13265 21635 13323 21641
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 17586 21672 17592 21684
rect 17547 21644 17592 21672
rect 17586 21632 17592 21644
rect 17644 21632 17650 21684
rect 4798 21604 4804 21616
rect 4448 21576 4804 21604
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4157 21539 4215 21545
rect 4157 21505 4169 21539
rect 4203 21505 4215 21539
rect 4157 21499 4215 21505
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 4080 21468 4108 21499
rect 4246 21496 4252 21548
rect 4304 21536 4310 21548
rect 4448 21545 4476 21576
rect 4798 21564 4804 21576
rect 4856 21604 4862 21616
rect 4856 21576 5856 21604
rect 4856 21564 4862 21576
rect 5828 21548 5856 21576
rect 4433 21539 4491 21545
rect 4304 21508 4349 21536
rect 4304 21496 4310 21508
rect 4433 21505 4445 21539
rect 4479 21505 4491 21539
rect 4433 21499 4491 21505
rect 5261 21539 5319 21545
rect 5261 21505 5273 21539
rect 5307 21505 5319 21539
rect 5261 21499 5319 21505
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21505 5411 21539
rect 5534 21536 5540 21548
rect 5495 21508 5540 21536
rect 5353 21499 5411 21505
rect 4522 21468 4528 21480
rect 2832 21440 2877 21468
rect 4080 21440 4528 21468
rect 2832 21428 2838 21440
rect 4522 21428 4528 21440
rect 4580 21428 4586 21480
rect 3237 21403 3295 21409
rect 3237 21369 3249 21403
rect 3283 21400 3295 21403
rect 3694 21400 3700 21412
rect 3283 21372 3700 21400
rect 3283 21369 3295 21372
rect 3237 21363 3295 21369
rect 3694 21360 3700 21372
rect 3752 21360 3758 21412
rect 3786 21332 3792 21344
rect 3747 21304 3792 21332
rect 3786 21292 3792 21304
rect 3844 21292 3850 21344
rect 5276 21332 5304 21499
rect 5368 21400 5396 21499
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 5718 21536 5724 21548
rect 5675 21508 5724 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 5718 21496 5724 21508
rect 5776 21496 5782 21548
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 7466 21536 7472 21548
rect 7524 21545 7530 21548
rect 7436 21508 7472 21536
rect 7466 21496 7472 21508
rect 7524 21499 7536 21545
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21536 7803 21539
rect 8205 21539 8263 21545
rect 8205 21536 8217 21539
rect 7791 21508 8217 21536
rect 7791 21505 7803 21508
rect 7745 21499 7803 21505
rect 8205 21505 8217 21508
rect 8251 21536 8263 21539
rect 8294 21536 8300 21548
rect 8251 21508 8300 21536
rect 8251 21505 8263 21508
rect 8205 21499 8263 21505
rect 7524 21496 7530 21499
rect 8294 21496 8300 21508
rect 8352 21496 8358 21548
rect 8478 21545 8484 21548
rect 8472 21499 8484 21545
rect 8536 21536 8542 21548
rect 10226 21536 10232 21548
rect 8536 21508 8572 21536
rect 10187 21508 10232 21536
rect 8478 21496 8484 21499
rect 8536 21496 8542 21508
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 11517 21539 11575 21545
rect 11517 21505 11529 21539
rect 11563 21536 11575 21539
rect 11882 21536 11888 21548
rect 11563 21508 11888 21536
rect 11563 21505 11575 21508
rect 11517 21499 11575 21505
rect 11882 21496 11888 21508
rect 11940 21496 11946 21548
rect 13446 21536 13452 21548
rect 13407 21508 13452 21536
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 16942 21536 16948 21548
rect 16903 21508 16948 21536
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 17770 21536 17776 21548
rect 17731 21508 17776 21536
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 10045 21471 10103 21477
rect 10045 21468 10057 21471
rect 9732 21440 10057 21468
rect 9732 21428 9738 21440
rect 10045 21437 10057 21440
rect 10091 21468 10103 21471
rect 10962 21468 10968 21480
rect 10091 21440 10968 21468
rect 10091 21437 10103 21440
rect 10045 21431 10103 21437
rect 10962 21428 10968 21440
rect 11020 21428 11026 21480
rect 6178 21400 6184 21412
rect 5368 21372 6184 21400
rect 6178 21360 6184 21372
rect 6236 21400 6242 21412
rect 6365 21403 6423 21409
rect 6365 21400 6377 21403
rect 6236 21372 6377 21400
rect 6236 21360 6242 21372
rect 6365 21369 6377 21372
rect 6411 21369 6423 21403
rect 6365 21363 6423 21369
rect 5626 21332 5632 21344
rect 5276 21304 5632 21332
rect 5626 21292 5632 21304
rect 5684 21292 5690 21344
rect 9582 21332 9588 21344
rect 9543 21304 9588 21332
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 11330 21292 11336 21344
rect 11388 21332 11394 21344
rect 11698 21332 11704 21344
rect 11388 21304 11704 21332
rect 11388 21292 11394 21304
rect 11698 21292 11704 21304
rect 11756 21292 11762 21344
rect 1104 21242 18860 21264
rect 1104 21190 3915 21242
rect 3967 21190 3979 21242
rect 4031 21190 4043 21242
rect 4095 21190 4107 21242
rect 4159 21190 4171 21242
rect 4223 21190 9846 21242
rect 9898 21190 9910 21242
rect 9962 21190 9974 21242
rect 10026 21190 10038 21242
rect 10090 21190 10102 21242
rect 10154 21190 15776 21242
rect 15828 21190 15840 21242
rect 15892 21190 15904 21242
rect 15956 21190 15968 21242
rect 16020 21190 16032 21242
rect 16084 21190 18860 21242
rect 1104 21168 18860 21190
rect 4522 21088 4528 21140
rect 4580 21128 4586 21140
rect 5261 21131 5319 21137
rect 5261 21128 5273 21131
rect 4580 21100 5273 21128
rect 4580 21088 4586 21100
rect 5261 21097 5273 21100
rect 5307 21097 5319 21131
rect 5261 21091 5319 21097
rect 16114 21088 16120 21140
rect 16172 21128 16178 21140
rect 17865 21131 17923 21137
rect 17865 21128 17877 21131
rect 16172 21100 17877 21128
rect 16172 21088 16178 21100
rect 17865 21097 17877 21100
rect 17911 21097 17923 21131
rect 17865 21091 17923 21097
rect 6178 20992 6184 21004
rect 6139 20964 6184 20992
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6454 20992 6460 21004
rect 6415 20964 6460 20992
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 11238 20952 11244 21004
rect 11296 20992 11302 21004
rect 11333 20995 11391 21001
rect 11333 20992 11345 20995
rect 11296 20964 11345 20992
rect 11296 20952 11302 20964
rect 11333 20961 11345 20964
rect 11379 20961 11391 20995
rect 11333 20955 11391 20961
rect 3881 20927 3939 20933
rect 3881 20893 3893 20927
rect 3927 20924 3939 20927
rect 4430 20924 4436 20936
rect 3927 20896 4436 20924
rect 3927 20893 3939 20896
rect 3881 20887 3939 20893
rect 4430 20884 4436 20896
rect 4488 20884 4494 20936
rect 7374 20884 7380 20936
rect 7432 20924 7438 20936
rect 7837 20927 7895 20933
rect 7837 20924 7849 20927
rect 7432 20896 7849 20924
rect 7432 20884 7438 20896
rect 7837 20893 7849 20896
rect 7883 20893 7895 20927
rect 8110 20924 8116 20936
rect 8071 20896 8116 20924
rect 7837 20887 7895 20893
rect 8110 20884 8116 20896
rect 8168 20884 8174 20936
rect 8294 20884 8300 20936
rect 8352 20924 8358 20936
rect 11606 20933 11612 20936
rect 10873 20927 10931 20933
rect 10873 20924 10885 20927
rect 8352 20896 10885 20924
rect 8352 20884 8358 20896
rect 10873 20893 10885 20896
rect 10919 20893 10931 20927
rect 10873 20887 10931 20893
rect 11600 20887 11612 20933
rect 11664 20924 11670 20936
rect 11664 20896 11700 20924
rect 11606 20884 11612 20887
rect 11664 20884 11670 20896
rect 12710 20884 12716 20936
rect 12768 20924 12774 20936
rect 13265 20927 13323 20933
rect 13265 20924 13277 20927
rect 12768 20896 13277 20924
rect 12768 20884 12774 20896
rect 13265 20893 13277 20896
rect 13311 20893 13323 20927
rect 13265 20887 13323 20893
rect 13354 20884 13360 20936
rect 13412 20924 13418 20936
rect 18049 20927 18107 20933
rect 18049 20924 18061 20927
rect 13412 20896 18061 20924
rect 13412 20884 13418 20896
rect 18049 20893 18061 20896
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 3786 20816 3792 20868
rect 3844 20856 3850 20868
rect 4126 20859 4184 20865
rect 4126 20856 4138 20859
rect 3844 20828 4138 20856
rect 3844 20816 3850 20828
rect 4126 20825 4138 20828
rect 4172 20825 4184 20859
rect 4126 20819 4184 20825
rect 8021 20859 8079 20865
rect 8021 20825 8033 20859
rect 8067 20856 8079 20859
rect 9582 20856 9588 20868
rect 8067 20828 9588 20856
rect 8067 20825 8079 20828
rect 8021 20819 8079 20825
rect 9582 20816 9588 20828
rect 9640 20816 9646 20868
rect 10628 20859 10686 20865
rect 10628 20825 10640 20859
rect 10674 20856 10686 20859
rect 10778 20856 10784 20868
rect 10674 20828 10784 20856
rect 10674 20825 10686 20828
rect 10628 20819 10686 20825
rect 10778 20816 10784 20828
rect 10836 20816 10842 20868
rect 7650 20788 7656 20800
rect 7611 20760 7656 20788
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 9490 20788 9496 20800
rect 9451 20760 9496 20788
rect 9490 20748 9496 20760
rect 9548 20748 9554 20800
rect 12713 20791 12771 20797
rect 12713 20757 12725 20791
rect 12759 20788 12771 20791
rect 13170 20788 13176 20800
rect 12759 20760 13176 20788
rect 12759 20757 12771 20760
rect 12713 20751 12771 20757
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 1104 20698 18860 20720
rect 1104 20646 6880 20698
rect 6932 20646 6944 20698
rect 6996 20646 7008 20698
rect 7060 20646 7072 20698
rect 7124 20646 7136 20698
rect 7188 20646 12811 20698
rect 12863 20646 12875 20698
rect 12927 20646 12939 20698
rect 12991 20646 13003 20698
rect 13055 20646 13067 20698
rect 13119 20646 18860 20698
rect 1104 20624 18860 20646
rect 3881 20587 3939 20593
rect 3881 20553 3893 20587
rect 3927 20584 3939 20587
rect 4246 20584 4252 20596
rect 3927 20556 4252 20584
rect 3927 20553 3939 20556
rect 3881 20547 3939 20553
rect 4246 20544 4252 20556
rect 4304 20544 4310 20596
rect 5721 20587 5779 20593
rect 5721 20553 5733 20587
rect 5767 20584 5779 20587
rect 7466 20584 7472 20596
rect 5767 20556 7472 20584
rect 5767 20553 5779 20556
rect 5721 20547 5779 20553
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 7745 20587 7803 20593
rect 7745 20553 7757 20587
rect 7791 20584 7803 20587
rect 8386 20584 8392 20596
rect 7791 20556 8392 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 8386 20544 8392 20556
rect 8444 20584 8450 20596
rect 8570 20584 8576 20596
rect 8444 20556 8576 20584
rect 8444 20544 8450 20556
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 10071 20587 10129 20593
rect 10071 20553 10083 20587
rect 10117 20584 10129 20587
rect 10226 20584 10232 20596
rect 10117 20556 10232 20584
rect 10117 20553 10129 20556
rect 10071 20547 10129 20553
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11422 20584 11428 20596
rect 11011 20556 11428 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 11422 20544 11428 20556
rect 11480 20544 11486 20596
rect 3602 20476 3608 20528
rect 3660 20516 3666 20528
rect 7561 20519 7619 20525
rect 3660 20488 3924 20516
rect 3660 20476 3666 20488
rect 3694 20448 3700 20460
rect 3655 20420 3700 20448
rect 3694 20408 3700 20420
rect 3752 20408 3758 20460
rect 3896 20457 3924 20488
rect 7561 20485 7573 20519
rect 7607 20516 7619 20519
rect 7650 20516 7656 20528
rect 7607 20488 7656 20516
rect 7607 20485 7619 20488
rect 7561 20479 7619 20485
rect 7650 20476 7656 20488
rect 7708 20476 7714 20528
rect 9490 20476 9496 20528
rect 9548 20516 9554 20528
rect 9861 20519 9919 20525
rect 9861 20516 9873 20519
rect 9548 20488 9873 20516
rect 9548 20476 9554 20488
rect 9861 20485 9873 20488
rect 9907 20485 9919 20519
rect 10244 20516 10272 20544
rect 10244 20488 10824 20516
rect 9861 20479 9919 20485
rect 3881 20451 3939 20457
rect 3881 20417 3893 20451
rect 3927 20417 3939 20451
rect 3881 20411 3939 20417
rect 5629 20451 5687 20457
rect 5629 20417 5641 20451
rect 5675 20448 5687 20451
rect 5718 20448 5724 20460
rect 5675 20420 5724 20448
rect 5675 20417 5687 20420
rect 5629 20411 5687 20417
rect 5718 20408 5724 20420
rect 5776 20408 5782 20460
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 6454 20448 6460 20460
rect 5859 20420 6460 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 6454 20408 6460 20420
rect 6512 20408 6518 20460
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20448 6699 20451
rect 7374 20448 7380 20460
rect 6687 20420 7380 20448
rect 6687 20417 6699 20420
rect 6641 20411 6699 20417
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 7834 20408 7840 20460
rect 7892 20448 7898 20460
rect 9030 20448 9036 20460
rect 7892 20420 7937 20448
rect 8991 20420 9036 20448
rect 7892 20408 7898 20420
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 10796 20457 10824 20488
rect 11882 20476 11888 20528
rect 11940 20516 11946 20528
rect 11977 20519 12035 20525
rect 11977 20516 11989 20519
rect 11940 20488 11989 20516
rect 11940 20476 11946 20488
rect 11977 20485 11989 20488
rect 12023 20516 12035 20519
rect 13081 20519 13139 20525
rect 13081 20516 13093 20519
rect 12023 20488 13093 20516
rect 12023 20485 12035 20488
rect 11977 20479 12035 20485
rect 13081 20485 13093 20488
rect 13127 20516 13139 20519
rect 15286 20516 15292 20528
rect 13127 20488 15292 20516
rect 13127 20485 13139 20488
rect 13081 20479 13139 20485
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 10689 20451 10747 20457
rect 10689 20448 10701 20451
rect 10060 20420 10701 20448
rect 7561 20315 7619 20321
rect 7561 20281 7573 20315
rect 7607 20312 7619 20315
rect 8478 20312 8484 20324
rect 7607 20284 8484 20312
rect 7607 20281 7619 20284
rect 7561 20275 7619 20281
rect 8478 20272 8484 20284
rect 8536 20272 8542 20324
rect 5994 20204 6000 20256
rect 6052 20244 6058 20256
rect 6457 20247 6515 20253
rect 6457 20244 6469 20247
rect 6052 20216 6469 20244
rect 6052 20204 6058 20216
rect 6457 20213 6469 20216
rect 6503 20213 6515 20247
rect 6457 20207 6515 20213
rect 8570 20204 8576 20256
rect 8628 20244 8634 20256
rect 8941 20247 8999 20253
rect 8941 20244 8953 20247
rect 8628 20216 8953 20244
rect 8628 20204 8634 20216
rect 8941 20213 8953 20216
rect 8987 20213 8999 20247
rect 8941 20207 8999 20213
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 10060 20253 10088 20420
rect 10689 20417 10701 20420
rect 10735 20417 10747 20451
rect 10689 20411 10747 20417
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20417 10839 20451
rect 10781 20411 10839 20417
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 12897 20451 12955 20457
rect 12897 20448 12909 20451
rect 12768 20420 12909 20448
rect 12768 20408 12774 20420
rect 12897 20417 12909 20420
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11330 20380 11336 20392
rect 11011 20352 11336 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 11330 20340 11336 20352
rect 11388 20340 11394 20392
rect 12158 20312 12164 20324
rect 12119 20284 12164 20312
rect 12158 20272 12164 20284
rect 12216 20272 12222 20324
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 9732 20216 10057 20244
rect 9732 20204 9738 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 10226 20204 10232 20256
rect 10284 20244 10290 20256
rect 10962 20244 10968 20256
rect 10284 20216 10968 20244
rect 10284 20204 10290 20216
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 1104 20154 18860 20176
rect 1104 20102 3915 20154
rect 3967 20102 3979 20154
rect 4031 20102 4043 20154
rect 4095 20102 4107 20154
rect 4159 20102 4171 20154
rect 4223 20102 9846 20154
rect 9898 20102 9910 20154
rect 9962 20102 9974 20154
rect 10026 20102 10038 20154
rect 10090 20102 10102 20154
rect 10154 20102 15776 20154
rect 15828 20102 15840 20154
rect 15892 20102 15904 20154
rect 15956 20102 15968 20154
rect 16020 20102 16032 20154
rect 16084 20102 18860 20154
rect 1104 20080 18860 20102
rect 7834 20000 7840 20052
rect 7892 20040 7898 20052
rect 8113 20043 8171 20049
rect 8113 20040 8125 20043
rect 7892 20012 8125 20040
rect 7892 20000 7898 20012
rect 8113 20009 8125 20012
rect 8159 20009 8171 20043
rect 10778 20040 10784 20052
rect 10739 20012 10784 20040
rect 8113 20003 8171 20009
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 10137 19975 10195 19981
rect 10137 19941 10149 19975
rect 10183 19972 10195 19975
rect 10686 19972 10692 19984
rect 10183 19944 10692 19972
rect 10183 19941 10195 19944
rect 10137 19935 10195 19941
rect 10686 19932 10692 19944
rect 10744 19932 10750 19984
rect 14737 19975 14795 19981
rect 14737 19941 14749 19975
rect 14783 19972 14795 19975
rect 15010 19972 15016 19984
rect 14783 19944 15016 19972
rect 14783 19941 14795 19944
rect 14737 19935 14795 19941
rect 15010 19932 15016 19944
rect 15068 19932 15074 19984
rect 10321 19907 10379 19913
rect 10321 19873 10333 19907
rect 10367 19904 10379 19907
rect 11330 19904 11336 19916
rect 10367 19876 11336 19904
rect 10367 19873 10379 19876
rect 10321 19867 10379 19873
rect 11330 19864 11336 19876
rect 11388 19864 11394 19916
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 8168 19808 8217 19836
rect 8168 19796 8174 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 9490 19796 9496 19848
rect 9548 19836 9554 19848
rect 9585 19839 9643 19845
rect 9585 19836 9597 19839
rect 9548 19808 9597 19836
rect 9548 19796 9554 19808
rect 9585 19805 9597 19808
rect 9631 19836 9643 19839
rect 10045 19839 10103 19845
rect 10045 19836 10057 19839
rect 9631 19808 10057 19836
rect 9631 19805 9643 19808
rect 9585 19799 9643 19805
rect 10045 19805 10057 19808
rect 10091 19805 10103 19839
rect 10781 19839 10839 19845
rect 10781 19836 10793 19839
rect 10045 19799 10103 19805
rect 10336 19808 10793 19836
rect 10336 19777 10364 19808
rect 10781 19805 10793 19808
rect 10827 19805 10839 19839
rect 10962 19836 10968 19848
rect 10923 19808 10968 19836
rect 10781 19799 10839 19805
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 15102 19796 15108 19848
rect 15160 19836 15166 19848
rect 15565 19839 15623 19845
rect 15565 19836 15577 19839
rect 15160 19808 15577 19836
rect 15160 19796 15166 19808
rect 15565 19805 15577 19808
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 15712 19808 15761 19836
rect 15712 19796 15718 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 10321 19771 10379 19777
rect 10321 19737 10333 19771
rect 10367 19737 10379 19771
rect 10321 19731 10379 19737
rect 12710 19728 12716 19780
rect 12768 19768 12774 19780
rect 14553 19771 14611 19777
rect 14553 19768 14565 19771
rect 12768 19740 14565 19768
rect 12768 19728 12774 19740
rect 14553 19737 14565 19740
rect 14599 19737 14611 19771
rect 14553 19731 14611 19737
rect 9490 19700 9496 19712
rect 9451 19672 9496 19700
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 15933 19703 15991 19709
rect 15933 19669 15945 19703
rect 15979 19700 15991 19703
rect 16666 19700 16672 19712
rect 15979 19672 16672 19700
rect 15979 19669 15991 19672
rect 15933 19663 15991 19669
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 1104 19610 18860 19632
rect 1104 19558 6880 19610
rect 6932 19558 6944 19610
rect 6996 19558 7008 19610
rect 7060 19558 7072 19610
rect 7124 19558 7136 19610
rect 7188 19558 12811 19610
rect 12863 19558 12875 19610
rect 12927 19558 12939 19610
rect 12991 19558 13003 19610
rect 13055 19558 13067 19610
rect 13119 19558 18860 19610
rect 1104 19536 18860 19558
rect 14737 19499 14795 19505
rect 14737 19465 14749 19499
rect 14783 19496 14795 19499
rect 15194 19496 15200 19508
rect 14783 19468 15200 19496
rect 14783 19465 14795 19468
rect 14737 19459 14795 19465
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 9493 19431 9551 19437
rect 9493 19397 9505 19431
rect 9539 19428 9551 19431
rect 9766 19428 9772 19440
rect 9539 19400 9772 19428
rect 9539 19397 9551 19400
rect 9493 19391 9551 19397
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 14277 19431 14335 19437
rect 14277 19397 14289 19431
rect 14323 19428 14335 19431
rect 15102 19428 15108 19440
rect 14323 19400 15108 19428
rect 14323 19397 14335 19400
rect 14277 19391 14335 19397
rect 15102 19388 15108 19400
rect 15160 19388 15166 19440
rect 9585 19363 9643 19369
rect 9585 19329 9597 19363
rect 9631 19360 9643 19363
rect 9674 19360 9680 19372
rect 9631 19332 9680 19360
rect 9631 19329 9643 19332
rect 9585 19323 9643 19329
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 12710 19320 12716 19372
rect 12768 19360 12774 19372
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12768 19332 12909 19360
rect 12768 19320 12774 19332
rect 12897 19329 12909 19332
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 14553 19363 14611 19369
rect 14553 19329 14565 19363
rect 14599 19360 14611 19363
rect 14599 19332 14964 19360
rect 14599 19329 14611 19332
rect 14553 19323 14611 19329
rect 13081 19295 13139 19301
rect 13081 19261 13093 19295
rect 13127 19292 13139 19295
rect 13354 19292 13360 19304
rect 13127 19264 13360 19292
rect 13127 19261 13139 19264
rect 13081 19255 13139 19261
rect 13354 19252 13360 19264
rect 13412 19292 13418 19304
rect 14366 19292 14372 19304
rect 13412 19264 14372 19292
rect 13412 19252 13418 19264
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 13170 19116 13176 19168
rect 13228 19156 13234 19168
rect 14277 19159 14335 19165
rect 14277 19156 14289 19159
rect 13228 19128 14289 19156
rect 13228 19116 13234 19128
rect 14277 19125 14289 19128
rect 14323 19125 14335 19159
rect 14476 19156 14504 19323
rect 14936 19224 14964 19332
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 16666 19360 16672 19372
rect 15068 19332 15240 19360
rect 16627 19332 16672 19360
rect 15068 19320 15074 19332
rect 15212 19301 15240 19332
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 15197 19295 15255 19301
rect 15197 19261 15209 19295
rect 15243 19261 15255 19295
rect 15197 19255 15255 19261
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 16206 19292 16212 19304
rect 15519 19264 16212 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 15378 19224 15384 19236
rect 14936 19196 15384 19224
rect 15378 19184 15384 19196
rect 15436 19184 15442 19236
rect 16114 19156 16120 19168
rect 14476 19128 16120 19156
rect 14277 19119 14335 19125
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 16850 19156 16856 19168
rect 16811 19128 16856 19156
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 1104 19066 18860 19088
rect 1104 19014 3915 19066
rect 3967 19014 3979 19066
rect 4031 19014 4043 19066
rect 4095 19014 4107 19066
rect 4159 19014 4171 19066
rect 4223 19014 9846 19066
rect 9898 19014 9910 19066
rect 9962 19014 9974 19066
rect 10026 19014 10038 19066
rect 10090 19014 10102 19066
rect 10154 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 15904 19066
rect 15956 19014 15968 19066
rect 16020 19014 16032 19066
rect 16084 19014 18860 19066
rect 1104 18992 18860 19014
rect 5626 18952 5632 18964
rect 5587 18924 5632 18952
rect 5626 18912 5632 18924
rect 5684 18912 5690 18964
rect 14369 18955 14427 18961
rect 14369 18921 14381 18955
rect 14415 18952 14427 18955
rect 15102 18952 15108 18964
rect 14415 18924 15108 18952
rect 14415 18921 14427 18924
rect 14369 18915 14427 18921
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 16209 18955 16267 18961
rect 16209 18952 16221 18955
rect 16172 18924 16221 18952
rect 16172 18912 16178 18924
rect 16209 18921 16221 18924
rect 16255 18921 16267 18955
rect 16209 18915 16267 18921
rect 12437 18887 12495 18893
rect 12437 18853 12449 18887
rect 12483 18884 12495 18887
rect 12526 18884 12532 18896
rect 12483 18856 12532 18884
rect 12483 18853 12495 18856
rect 12437 18847 12495 18853
rect 12526 18844 12532 18856
rect 12584 18844 12590 18896
rect 13170 18816 13176 18828
rect 13131 18788 13176 18816
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 5718 18748 5724 18760
rect 5679 18720 5724 18748
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 12066 18708 12072 18760
rect 12124 18748 12130 18760
rect 12253 18751 12311 18757
rect 12253 18748 12265 18751
rect 12124 18720 12265 18748
rect 12124 18708 12130 18720
rect 12253 18717 12265 18720
rect 12299 18717 12311 18751
rect 12434 18748 12440 18760
rect 12395 18720 12440 18748
rect 12253 18711 12311 18717
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 13354 18748 13360 18760
rect 13315 18720 13360 18748
rect 13354 18708 13360 18720
rect 13412 18708 13418 18760
rect 14918 18708 14924 18760
rect 14976 18748 14982 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 14976 18720 15761 18748
rect 14976 18708 14982 18720
rect 15749 18717 15761 18720
rect 15795 18748 15807 18751
rect 16758 18748 16764 18760
rect 15795 18720 16764 18748
rect 15795 18717 15807 18720
rect 15749 18711 15807 18717
rect 16758 18708 16764 18720
rect 16816 18748 16822 18760
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 16816 18720 17601 18748
rect 16816 18708 16822 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 15470 18680 15476 18692
rect 15528 18689 15534 18692
rect 15440 18652 15476 18680
rect 15470 18640 15476 18652
rect 15528 18643 15540 18689
rect 15528 18640 15534 18643
rect 16850 18640 16856 18692
rect 16908 18680 16914 18692
rect 17322 18683 17380 18689
rect 17322 18680 17334 18683
rect 16908 18652 17334 18680
rect 16908 18640 16914 18652
rect 17322 18649 17334 18652
rect 17368 18649 17380 18683
rect 17322 18643 17380 18649
rect 13354 18572 13360 18624
rect 13412 18612 13418 18624
rect 13541 18615 13599 18621
rect 13541 18612 13553 18615
rect 13412 18584 13553 18612
rect 13412 18572 13418 18584
rect 13541 18581 13553 18584
rect 13587 18581 13599 18615
rect 13541 18575 13599 18581
rect 1104 18522 18860 18544
rect 1104 18470 6880 18522
rect 6932 18470 6944 18522
rect 6996 18470 7008 18522
rect 7060 18470 7072 18522
rect 7124 18470 7136 18522
rect 7188 18470 12811 18522
rect 12863 18470 12875 18522
rect 12927 18470 12939 18522
rect 12991 18470 13003 18522
rect 13055 18470 13067 18522
rect 13119 18470 18860 18522
rect 1104 18448 18860 18470
rect 4893 18411 4951 18417
rect 4893 18377 4905 18411
rect 4939 18408 4951 18411
rect 5534 18408 5540 18420
rect 4939 18380 5540 18408
rect 4939 18377 4951 18380
rect 4893 18371 4951 18377
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 8202 18408 8208 18420
rect 5736 18380 8208 18408
rect 4246 18232 4252 18284
rect 4304 18272 4310 18284
rect 4801 18275 4859 18281
rect 4801 18272 4813 18275
rect 4304 18244 4813 18272
rect 4304 18232 4310 18244
rect 4801 18241 4813 18244
rect 4847 18272 4859 18275
rect 5258 18272 5264 18284
rect 4847 18244 5264 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5736 18281 5764 18380
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 6362 18300 6368 18352
rect 6420 18340 6426 18352
rect 7469 18343 7527 18349
rect 7469 18340 7481 18343
rect 6420 18312 7481 18340
rect 6420 18300 6426 18312
rect 7469 18309 7481 18312
rect 7515 18309 7527 18343
rect 7469 18303 7527 18309
rect 14090 18300 14096 18352
rect 14148 18340 14154 18352
rect 14148 18312 14780 18340
rect 14148 18300 14154 18312
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18241 5779 18275
rect 5721 18235 5779 18241
rect 6457 18275 6515 18281
rect 6457 18241 6469 18275
rect 6503 18241 6515 18275
rect 6457 18235 6515 18241
rect 1394 18068 1400 18080
rect 1355 18040 1400 18068
rect 1394 18028 1400 18040
rect 1452 18028 1458 18080
rect 5534 18068 5540 18080
rect 5495 18040 5540 18068
rect 5534 18028 5540 18040
rect 5592 18068 5598 18080
rect 5810 18068 5816 18080
rect 5592 18040 5816 18068
rect 5592 18028 5598 18040
rect 5810 18028 5816 18040
rect 5868 18028 5874 18080
rect 6472 18068 6500 18235
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 6604 18244 6649 18272
rect 6604 18232 6610 18244
rect 6730 18232 6736 18284
rect 6788 18272 6794 18284
rect 7193 18275 7251 18281
rect 6788 18244 6833 18272
rect 6788 18232 6794 18244
rect 7193 18241 7205 18275
rect 7239 18241 7251 18275
rect 12434 18272 12440 18284
rect 12395 18244 12440 18272
rect 7193 18235 7251 18241
rect 7208 18204 7236 18235
rect 12434 18232 12440 18244
rect 12492 18232 12498 18284
rect 14642 18272 14648 18284
rect 14700 18281 14706 18284
rect 14612 18244 14648 18272
rect 14642 18232 14648 18244
rect 14700 18235 14712 18281
rect 14752 18272 14780 18312
rect 15194 18300 15200 18352
rect 15252 18340 15258 18352
rect 15252 18312 15792 18340
rect 15252 18300 15258 18312
rect 14918 18272 14924 18284
rect 14752 18244 14924 18272
rect 14700 18232 14706 18235
rect 14918 18232 14924 18244
rect 14976 18232 14982 18284
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15764 18281 15792 18312
rect 15381 18275 15439 18281
rect 15381 18272 15393 18275
rect 15344 18244 15393 18272
rect 15344 18232 15350 18244
rect 15381 18241 15393 18244
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18241 15715 18275
rect 15657 18235 15715 18241
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 6748 18176 7236 18204
rect 7469 18207 7527 18213
rect 6748 18145 6776 18176
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7650 18204 7656 18216
rect 7515 18176 7656 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12621 18207 12679 18213
rect 12621 18204 12633 18207
rect 12124 18176 12633 18204
rect 12124 18164 12130 18176
rect 12621 18173 12633 18176
rect 12667 18173 12679 18207
rect 15580 18204 15608 18235
rect 12621 18167 12679 18173
rect 15120 18176 15608 18204
rect 6733 18139 6791 18145
rect 6733 18105 6745 18139
rect 6779 18105 6791 18139
rect 7190 18136 7196 18148
rect 6733 18099 6791 18105
rect 6840 18108 7196 18136
rect 6840 18068 6868 18108
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 6472 18040 6868 18068
rect 6914 18028 6920 18080
rect 6972 18068 6978 18080
rect 7285 18071 7343 18077
rect 7285 18068 7297 18071
rect 6972 18040 7297 18068
rect 6972 18028 6978 18040
rect 7285 18037 7297 18040
rect 7331 18037 7343 18071
rect 12250 18068 12256 18080
rect 12211 18040 12256 18068
rect 7285 18031 7343 18037
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 13541 18071 13599 18077
rect 13541 18037 13553 18071
rect 13587 18068 13599 18071
rect 14550 18068 14556 18080
rect 13587 18040 14556 18068
rect 13587 18037 13599 18040
rect 13541 18031 13599 18037
rect 14550 18028 14556 18040
rect 14608 18068 14614 18080
rect 15120 18068 15148 18176
rect 15672 18136 15700 18235
rect 16206 18232 16212 18284
rect 16264 18272 16270 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16264 18244 16865 18272
rect 16264 18232 16270 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 16298 18164 16304 18216
rect 16356 18204 16362 18216
rect 17037 18207 17095 18213
rect 17037 18204 17049 18207
rect 16356 18176 17049 18204
rect 16356 18164 16362 18176
rect 17037 18173 17049 18176
rect 17083 18173 17095 18207
rect 17037 18167 17095 18173
rect 17402 18136 17408 18148
rect 15672 18108 17408 18136
rect 17402 18096 17408 18108
rect 17460 18096 17466 18148
rect 14608 18040 15148 18068
rect 14608 18028 14614 18040
rect 15194 18028 15200 18080
rect 15252 18068 15258 18080
rect 16025 18071 16083 18077
rect 16025 18068 16037 18071
rect 15252 18040 16037 18068
rect 15252 18028 15258 18040
rect 16025 18037 16037 18040
rect 16071 18037 16083 18071
rect 16666 18068 16672 18080
rect 16627 18040 16672 18068
rect 16025 18031 16083 18037
rect 16666 18028 16672 18040
rect 16724 18028 16730 18080
rect 1104 17978 18860 18000
rect 1104 17926 3915 17978
rect 3967 17926 3979 17978
rect 4031 17926 4043 17978
rect 4095 17926 4107 17978
rect 4159 17926 4171 17978
rect 4223 17926 9846 17978
rect 9898 17926 9910 17978
rect 9962 17926 9974 17978
rect 10026 17926 10038 17978
rect 10090 17926 10102 17978
rect 10154 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 15904 17978
rect 15956 17926 15968 17978
rect 16020 17926 16032 17978
rect 16084 17926 18860 17978
rect 1104 17904 18860 17926
rect 4890 17824 4896 17876
rect 4948 17864 4954 17876
rect 4985 17867 5043 17873
rect 4985 17864 4997 17867
rect 4948 17836 4997 17864
rect 4948 17824 4954 17836
rect 4985 17833 4997 17836
rect 5031 17833 5043 17867
rect 7190 17864 7196 17876
rect 7151 17836 7196 17864
rect 4985 17827 5043 17833
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 11514 17864 11520 17876
rect 10827 17836 11520 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 4433 17799 4491 17805
rect 4433 17765 4445 17799
rect 4479 17796 4491 17799
rect 4614 17796 4620 17808
rect 4479 17768 4620 17796
rect 4479 17765 4491 17768
rect 4433 17759 4491 17765
rect 4614 17756 4620 17768
rect 4672 17756 4678 17808
rect 5902 17756 5908 17808
rect 5960 17796 5966 17808
rect 9674 17796 9680 17808
rect 5960 17768 9680 17796
rect 5960 17756 5966 17768
rect 9674 17756 9680 17768
rect 9732 17796 9738 17808
rect 10502 17796 10508 17808
rect 9732 17768 10508 17796
rect 9732 17756 9738 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 6178 17728 6184 17740
rect 6091 17700 6184 17728
rect 6178 17688 6184 17700
rect 6236 17728 6242 17740
rect 6730 17728 6736 17740
rect 6236 17700 6736 17728
rect 6236 17688 6242 17700
rect 6730 17688 6736 17700
rect 6788 17688 6794 17740
rect 7558 17688 7564 17740
rect 7616 17728 7622 17740
rect 8021 17731 8079 17737
rect 8021 17728 8033 17731
rect 7616 17700 8033 17728
rect 7616 17688 7622 17700
rect 8021 17697 8033 17700
rect 8067 17697 8079 17731
rect 10796 17728 10824 17827
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 12618 17864 12624 17876
rect 11624 17836 12624 17864
rect 11624 17728 11652 17836
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 15102 17824 15108 17876
rect 15160 17864 15166 17876
rect 16117 17867 16175 17873
rect 16117 17864 16129 17867
rect 15160 17836 16129 17864
rect 15160 17824 15166 17836
rect 16117 17833 16129 17836
rect 16163 17833 16175 17867
rect 16117 17827 16175 17833
rect 11790 17756 11796 17808
rect 11848 17796 11854 17808
rect 11977 17799 12035 17805
rect 11977 17796 11989 17799
rect 11848 17768 11989 17796
rect 11848 17756 11854 17768
rect 11977 17765 11989 17768
rect 12023 17765 12035 17799
rect 11977 17759 12035 17765
rect 12710 17756 12716 17808
rect 12768 17756 12774 17808
rect 15378 17756 15384 17808
rect 15436 17796 15442 17808
rect 15473 17799 15531 17805
rect 15473 17796 15485 17799
rect 15436 17768 15485 17796
rect 15436 17756 15442 17768
rect 15473 17765 15485 17768
rect 15519 17765 15531 17799
rect 15473 17759 15531 17765
rect 8021 17691 8079 17697
rect 9048 17700 10824 17728
rect 11247 17700 11652 17728
rect 12069 17731 12127 17737
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4706 17660 4712 17672
rect 4295 17632 4712 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4706 17620 4712 17632
rect 4764 17660 4770 17672
rect 5166 17660 5172 17672
rect 4764 17632 5172 17660
rect 4764 17620 4770 17632
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6270 17660 6276 17672
rect 6231 17632 6276 17660
rect 6270 17620 6276 17632
rect 6328 17620 6334 17672
rect 6454 17660 6460 17672
rect 6415 17632 6460 17660
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 8202 17660 8208 17672
rect 8115 17632 8208 17660
rect 8202 17620 8208 17632
rect 8260 17660 8266 17672
rect 9048 17660 9076 17700
rect 8260 17632 9076 17660
rect 8260 17620 8266 17632
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9732 17632 9781 17660
rect 9732 17620 9738 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 10962 17660 10968 17672
rect 9999 17632 10968 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 7374 17592 7380 17604
rect 7335 17564 7380 17592
rect 7374 17552 7380 17564
rect 7432 17552 7438 17604
rect 7561 17595 7619 17601
rect 7561 17561 7573 17595
rect 7607 17592 7619 17595
rect 7742 17592 7748 17604
rect 7607 17564 7748 17592
rect 7607 17561 7619 17564
rect 7561 17555 7619 17561
rect 7742 17552 7748 17564
rect 7800 17592 7806 17604
rect 10873 17595 10931 17601
rect 7800 17564 9996 17592
rect 7800 17552 7806 17564
rect 6638 17524 6644 17536
rect 6599 17496 6644 17524
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 9858 17524 9864 17536
rect 9819 17496 9864 17524
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 9968 17524 9996 17564
rect 10873 17561 10885 17595
rect 10919 17592 10931 17595
rect 11146 17592 11152 17604
rect 10919 17564 11152 17592
rect 10919 17561 10931 17564
rect 10873 17555 10931 17561
rect 11146 17552 11152 17564
rect 11204 17552 11210 17604
rect 11247 17524 11275 17700
rect 12069 17697 12081 17731
rect 12115 17728 12127 17731
rect 12250 17728 12256 17740
rect 12115 17700 12256 17728
rect 12115 17697 12127 17700
rect 12069 17691 12127 17697
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 11698 17660 11704 17672
rect 11659 17632 11704 17660
rect 11698 17620 11704 17632
rect 11756 17620 11762 17672
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17629 11851 17663
rect 12526 17660 12532 17672
rect 11793 17623 11851 17629
rect 12176 17632 12532 17660
rect 11808 17592 11836 17623
rect 12176 17592 12204 17632
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 12728 17669 12756 17756
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17629 12771 17663
rect 12713 17623 12771 17629
rect 11808 17564 12204 17592
rect 12342 17552 12348 17604
rect 12400 17592 12406 17604
rect 12728 17592 12756 17623
rect 12802 17620 12808 17672
rect 12860 17660 12866 17672
rect 13354 17660 13360 17672
rect 12860 17632 12905 17660
rect 13315 17632 13360 17660
rect 12860 17620 12866 17632
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 14090 17660 14096 17672
rect 14051 17632 14096 17660
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14338 17595 14396 17601
rect 14338 17592 14350 17595
rect 12400 17564 12756 17592
rect 13556 17564 14350 17592
rect 12400 17552 12406 17564
rect 11514 17524 11520 17536
rect 9968 17496 11275 17524
rect 11475 17496 11520 17524
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13556 17533 13584 17564
rect 14338 17561 14350 17564
rect 14384 17592 14396 17595
rect 14826 17592 14832 17604
rect 14384 17564 14832 17592
rect 14384 17561 14396 17564
rect 14338 17555 14396 17561
rect 14826 17552 14832 17564
rect 14884 17552 14890 17604
rect 15488 17592 15516 17759
rect 16206 17688 16212 17740
rect 16264 17728 16270 17740
rect 16390 17728 16396 17740
rect 16264 17700 16396 17728
rect 16264 17688 16270 17700
rect 16390 17688 16396 17700
rect 16448 17728 16454 17740
rect 16448 17700 16988 17728
rect 16448 17688 16454 17700
rect 16114 17620 16120 17672
rect 16172 17660 16178 17672
rect 16960 17669 16988 17700
rect 16761 17663 16819 17669
rect 16761 17660 16773 17663
rect 16172 17632 16773 17660
rect 16172 17620 16178 17632
rect 16761 17629 16773 17632
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17629 17003 17663
rect 16945 17623 17003 17629
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17660 17187 17663
rect 17773 17663 17831 17669
rect 17773 17660 17785 17663
rect 17175 17632 17785 17660
rect 17175 17629 17187 17632
rect 17129 17623 17187 17629
rect 17773 17629 17785 17632
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 16298 17592 16304 17604
rect 15488 17564 16304 17592
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 13541 17527 13599 17533
rect 13541 17493 13553 17527
rect 13587 17493 13599 17527
rect 15930 17524 15936 17536
rect 15891 17496 15936 17524
rect 13541 17487 13599 17493
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 16114 17533 16120 17536
rect 16101 17527 16120 17533
rect 16101 17493 16113 17527
rect 16101 17487 16120 17493
rect 16114 17484 16120 17487
rect 16172 17484 16178 17536
rect 17586 17524 17592 17536
rect 17547 17496 17592 17524
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 1104 17434 18860 17456
rect 1104 17382 6880 17434
rect 6932 17382 6944 17434
rect 6996 17382 7008 17434
rect 7060 17382 7072 17434
rect 7124 17382 7136 17434
rect 7188 17382 12811 17434
rect 12863 17382 12875 17434
rect 12927 17382 12939 17434
rect 12991 17382 13003 17434
rect 13055 17382 13067 17434
rect 13119 17382 18860 17434
rect 1104 17360 18860 17382
rect 4614 17320 4620 17332
rect 4264 17292 4620 17320
rect 4154 17184 4160 17196
rect 4115 17156 4160 17184
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4264 17193 4292 17292
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 5224 17292 11621 17320
rect 5224 17280 5230 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 14553 17323 14611 17329
rect 14553 17289 14565 17323
rect 14599 17320 14611 17323
rect 14642 17320 14648 17332
rect 14599 17292 14648 17320
rect 14599 17289 14611 17292
rect 14553 17283 14611 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 15528 17292 15577 17320
rect 15528 17280 15534 17292
rect 15565 17289 15577 17292
rect 15611 17289 15623 17323
rect 16666 17320 16672 17332
rect 15565 17283 15623 17289
rect 16546 17292 16672 17320
rect 5534 17252 5540 17264
rect 5000 17224 5540 17252
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17153 4307 17187
rect 4249 17147 4307 17153
rect 4341 17190 4399 17196
rect 4341 17156 4353 17190
rect 4387 17156 4399 17190
rect 4341 17150 4399 17156
rect 4525 17187 4583 17193
rect 4525 17153 4537 17187
rect 4571 17184 4583 17187
rect 5000 17184 5028 17224
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 6638 17261 6644 17264
rect 6632 17252 6644 17261
rect 6599 17224 6644 17252
rect 6632 17215 6644 17224
rect 6638 17212 6644 17215
rect 6696 17212 6702 17264
rect 10781 17255 10839 17261
rect 10781 17221 10793 17255
rect 10827 17252 10839 17255
rect 12342 17252 12348 17264
rect 10827 17224 12348 17252
rect 10827 17221 10839 17224
rect 10781 17215 10839 17221
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 15930 17252 15936 17264
rect 14660 17224 15936 17252
rect 5166 17184 5172 17196
rect 4571 17156 5028 17184
rect 5127 17156 5172 17184
rect 4571 17153 4583 17156
rect 3602 17076 3608 17128
rect 3660 17116 3666 17128
rect 4356 17116 4384 17150
rect 4525 17147 4583 17153
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5276 17156 5365 17184
rect 3660 17088 4384 17116
rect 3660 17076 3666 17088
rect 4614 17076 4620 17128
rect 4672 17116 4678 17128
rect 5276 17116 5304 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 8202 17184 8208 17196
rect 8163 17156 8208 17184
rect 5353 17147 5411 17153
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 8386 17184 8392 17196
rect 8347 17156 8392 17184
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 8570 17184 8576 17196
rect 8531 17156 8576 17184
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 8754 17184 8760 17196
rect 8715 17156 8760 17184
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 9858 17184 9864 17196
rect 9819 17156 9864 17184
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17184 10103 17187
rect 10226 17184 10232 17196
rect 10091 17156 10232 17184
rect 10091 17153 10103 17156
rect 10045 17147 10103 17153
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 11790 17184 11796 17196
rect 11624 17156 11796 17184
rect 5442 17116 5448 17128
rect 4672 17088 5304 17116
rect 5403 17088 5448 17116
rect 4672 17076 4678 17088
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 6365 17119 6423 17125
rect 6365 17085 6377 17119
rect 6411 17085 6423 17119
rect 6365 17079 6423 17085
rect 3786 17008 3792 17060
rect 3844 17048 3850 17060
rect 6380 17048 6408 17079
rect 7374 17076 7380 17128
rect 7432 17116 7438 17128
rect 8481 17119 8539 17125
rect 8481 17116 8493 17119
rect 7432 17088 8493 17116
rect 7432 17076 7438 17088
rect 8481 17085 8493 17088
rect 8527 17085 8539 17119
rect 8481 17079 8539 17085
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17116 10195 17119
rect 10686 17116 10692 17128
rect 10183 17088 10692 17116
rect 10183 17085 10195 17088
rect 10137 17079 10195 17085
rect 10686 17076 10692 17088
rect 10744 17076 10750 17128
rect 3844 17020 6408 17048
rect 3844 17008 3850 17020
rect 3881 16983 3939 16989
rect 3881 16949 3893 16983
rect 3927 16980 3939 16983
rect 4246 16980 4252 16992
rect 3927 16952 4252 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 4338 16940 4344 16992
rect 4396 16980 4402 16992
rect 4985 16983 5043 16989
rect 4985 16980 4997 16983
rect 4396 16952 4997 16980
rect 4396 16940 4402 16952
rect 4985 16949 4997 16952
rect 5031 16949 5043 16983
rect 6380 16980 6408 17020
rect 10965 17051 11023 17057
rect 10965 17017 10977 17051
rect 11011 17048 11023 17051
rect 11146 17048 11152 17060
rect 11011 17020 11152 17048
rect 11011 17017 11023 17020
rect 10965 17011 11023 17017
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 11624 17048 11652 17156
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17184 12219 17187
rect 12250 17184 12256 17196
rect 12207 17156 12256 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 11698 17076 11704 17128
rect 11756 17116 11762 17128
rect 11900 17116 11928 17147
rect 12250 17144 12256 17156
rect 12308 17144 12314 17196
rect 13446 17144 13452 17196
rect 13504 17184 13510 17196
rect 13725 17187 13783 17193
rect 13725 17184 13737 17187
rect 13504 17156 13737 17184
rect 13504 17144 13510 17156
rect 13725 17153 13737 17156
rect 13771 17153 13783 17187
rect 13725 17147 13783 17153
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 11756 17088 12633 17116
rect 11756 17076 11762 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 13262 17116 13268 17128
rect 13127 17088 13268 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 13262 17076 13268 17088
rect 13320 17116 13326 17128
rect 13541 17119 13599 17125
rect 13541 17116 13553 17119
rect 13320 17088 13553 17116
rect 13320 17076 13326 17088
rect 13541 17085 13553 17088
rect 13587 17085 13599 17119
rect 14660 17116 14688 17224
rect 15930 17212 15936 17224
rect 15988 17212 15994 17264
rect 14826 17184 14832 17196
rect 14787 17156 14832 17184
rect 14826 17144 14832 17156
rect 14884 17144 14890 17196
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17184 15071 17187
rect 15194 17184 15200 17196
rect 15059 17156 15200 17184
rect 15059 17153 15071 17156
rect 15013 17147 15071 17153
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17184 15807 17187
rect 16546 17184 16574 17292
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 17954 17280 17960 17332
rect 18012 17320 18018 17332
rect 18049 17323 18107 17329
rect 18049 17320 18061 17323
rect 18012 17292 18061 17320
rect 18012 17280 18018 17292
rect 18049 17289 18061 17292
rect 18095 17289 18107 17323
rect 18049 17283 18107 17289
rect 15795 17156 16574 17184
rect 16669 17187 16727 17193
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 16669 17153 16681 17187
rect 16715 17184 16727 17187
rect 16758 17184 16764 17196
rect 16715 17156 16764 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 16936 17187 16994 17193
rect 16936 17153 16948 17187
rect 16982 17184 16994 17187
rect 17310 17184 17316 17196
rect 16982 17156 17316 17184
rect 16982 17153 16994 17156
rect 16936 17147 16994 17153
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 14737 17119 14795 17125
rect 14737 17116 14749 17119
rect 14660 17088 14749 17116
rect 13541 17079 13599 17085
rect 14737 17085 14749 17088
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17116 14979 17119
rect 16022 17116 16028 17128
rect 14967 17088 16028 17116
rect 14967 17085 14979 17088
rect 14921 17079 14979 17085
rect 16022 17076 16028 17088
rect 16080 17076 16086 17128
rect 12250 17048 12256 17060
rect 11624 17020 12256 17048
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 12710 17048 12716 17060
rect 12671 17020 12716 17048
rect 12710 17008 12716 17020
rect 12768 17048 12774 17060
rect 13446 17048 13452 17060
rect 12768 17020 13452 17048
rect 12768 17008 12774 17020
rect 13446 17008 13452 17020
rect 13504 17008 13510 17060
rect 7006 16980 7012 16992
rect 6380 16952 7012 16980
rect 4985 16943 5043 16949
rect 7006 16940 7012 16952
rect 7064 16940 7070 16992
rect 7745 16983 7803 16989
rect 7745 16949 7757 16983
rect 7791 16980 7803 16983
rect 8018 16980 8024 16992
rect 7791 16952 8024 16980
rect 7791 16949 7803 16952
rect 7745 16943 7803 16949
rect 8018 16940 8024 16952
rect 8076 16940 8082 16992
rect 8938 16980 8944 16992
rect 8899 16952 8944 16980
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 9674 16980 9680 16992
rect 9635 16952 9680 16980
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 12069 16983 12127 16989
rect 12069 16949 12081 16983
rect 12115 16980 12127 16983
rect 12618 16980 12624 16992
rect 12115 16952 12624 16980
rect 12115 16949 12127 16952
rect 12069 16943 12127 16949
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 13909 16983 13967 16989
rect 13909 16949 13921 16983
rect 13955 16980 13967 16983
rect 15010 16980 15016 16992
rect 13955 16952 15016 16980
rect 13955 16949 13967 16952
rect 13909 16943 13967 16949
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 1104 16890 18860 16912
rect 1104 16838 3915 16890
rect 3967 16838 3979 16890
rect 4031 16838 4043 16890
rect 4095 16838 4107 16890
rect 4159 16838 4171 16890
rect 4223 16838 9846 16890
rect 9898 16838 9910 16890
rect 9962 16838 9974 16890
rect 10026 16838 10038 16890
rect 10090 16838 10102 16890
rect 10154 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 15904 16890
rect 15956 16838 15968 16890
rect 16020 16838 16032 16890
rect 16084 16838 18860 16890
rect 1104 16816 18860 16838
rect 3237 16779 3295 16785
rect 3237 16745 3249 16779
rect 3283 16776 3295 16779
rect 5166 16776 5172 16788
rect 3283 16748 5172 16776
rect 3283 16745 3295 16748
rect 3237 16739 3295 16745
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 8294 16776 8300 16788
rect 7064 16748 8300 16776
rect 7064 16736 7070 16748
rect 8294 16736 8300 16748
rect 8352 16776 8358 16788
rect 10686 16776 10692 16788
rect 8352 16748 9352 16776
rect 10647 16748 10692 16776
rect 8352 16736 8358 16748
rect 6270 16668 6276 16720
rect 6328 16668 6334 16720
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3510 16572 3516 16584
rect 3007 16544 3516 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3510 16532 3516 16544
rect 3568 16572 3574 16584
rect 3568 16544 3740 16572
rect 3568 16532 3574 16544
rect 3237 16507 3295 16513
rect 3237 16473 3249 16507
rect 3283 16504 3295 16507
rect 3326 16504 3332 16516
rect 3283 16476 3332 16504
rect 3283 16473 3295 16476
rect 3237 16467 3295 16473
rect 3326 16464 3332 16476
rect 3384 16464 3390 16516
rect 3712 16504 3740 16544
rect 3786 16532 3792 16584
rect 3844 16572 3850 16584
rect 4338 16581 4344 16584
rect 4065 16575 4123 16581
rect 4065 16572 4077 16575
rect 3844 16544 4077 16572
rect 3844 16532 3850 16544
rect 4065 16541 4077 16544
rect 4111 16541 4123 16575
rect 4332 16572 4344 16581
rect 4299 16544 4344 16572
rect 4065 16535 4123 16541
rect 4332 16535 4344 16544
rect 4338 16532 4344 16535
rect 4396 16532 4402 16584
rect 6288 16581 6316 16668
rect 9324 16652 9352 16748
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11238 16736 11244 16788
rect 11296 16776 11302 16788
rect 12342 16776 12348 16788
rect 11296 16748 12348 16776
rect 11296 16736 11302 16748
rect 12342 16736 12348 16748
rect 12400 16776 12406 16788
rect 14090 16776 14096 16788
rect 12400 16748 14096 16776
rect 12400 16736 12406 16748
rect 14090 16736 14096 16748
rect 14148 16776 14154 16788
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 14148 16748 14197 16776
rect 14148 16736 14154 16748
rect 14185 16745 14197 16748
rect 14231 16745 14243 16779
rect 14185 16739 14243 16745
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 16816 16748 17448 16776
rect 16816 16736 16822 16748
rect 12250 16668 12256 16720
rect 12308 16708 12314 16720
rect 13081 16711 13139 16717
rect 13081 16708 13093 16711
rect 12308 16680 13093 16708
rect 12308 16668 12314 16680
rect 13081 16677 13093 16680
rect 13127 16677 13139 16711
rect 13262 16708 13268 16720
rect 13223 16680 13268 16708
rect 13081 16671 13139 16677
rect 13262 16668 13268 16680
rect 13320 16668 13326 16720
rect 7006 16640 7012 16652
rect 6967 16612 7012 16640
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 9306 16640 9312 16652
rect 9219 16612 9312 16640
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 11238 16640 11244 16652
rect 11199 16612 11244 16640
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 13446 16600 13452 16652
rect 13504 16640 13510 16652
rect 17420 16649 17448 16748
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13504 16612 13553 16640
rect 13504 16600 13510 16612
rect 13541 16609 13553 16612
rect 13587 16609 13599 16643
rect 13541 16603 13599 16609
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16609 17463 16643
rect 17405 16603 17463 16609
rect 6181 16575 6239 16581
rect 6181 16572 6193 16575
rect 5828 16544 6193 16572
rect 4890 16504 4896 16516
rect 3712 16476 4896 16504
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 3053 16439 3111 16445
rect 3053 16405 3065 16439
rect 3099 16436 3111 16439
rect 4154 16436 4160 16448
rect 3099 16408 4160 16436
rect 3099 16405 3111 16408
rect 3053 16399 3111 16405
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 5445 16439 5503 16445
rect 5445 16405 5457 16439
rect 5491 16436 5503 16439
rect 5718 16436 5724 16448
rect 5491 16408 5724 16436
rect 5491 16405 5503 16408
rect 5445 16399 5503 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 5828 16436 5856 16544
rect 6181 16541 6193 16544
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16541 6331 16575
rect 6273 16535 6331 16541
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 6549 16575 6607 16581
rect 6420 16544 6465 16572
rect 6420 16532 6426 16544
rect 6549 16541 6561 16575
rect 6595 16572 6607 16575
rect 7558 16572 7564 16584
rect 6595 16544 7564 16572
rect 6595 16541 6607 16544
rect 6549 16535 6607 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 8754 16532 8760 16584
rect 8812 16572 8818 16584
rect 10134 16572 10140 16584
rect 8812 16544 10140 16572
rect 8812 16532 8818 16544
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 15010 16572 15016 16584
rect 14971 16544 15016 16572
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 17149 16575 17207 16581
rect 17149 16541 17161 16575
rect 17195 16572 17207 16575
rect 17586 16572 17592 16584
rect 17195 16544 17592 16572
rect 17195 16541 17207 16544
rect 17149 16535 17207 16541
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 5905 16507 5963 16513
rect 5905 16473 5917 16507
rect 5951 16504 5963 16507
rect 7254 16507 7312 16513
rect 7254 16504 7266 16507
rect 5951 16476 7266 16504
rect 5951 16473 5963 16476
rect 5905 16467 5963 16473
rect 7254 16473 7266 16476
rect 7300 16473 7312 16507
rect 7254 16467 7312 16473
rect 9576 16507 9634 16513
rect 9576 16473 9588 16507
rect 9622 16504 9634 16507
rect 9674 16504 9680 16516
rect 9622 16476 9680 16504
rect 9622 16473 9634 16476
rect 9576 16467 9634 16473
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 11508 16507 11566 16513
rect 11508 16473 11520 16507
rect 11554 16504 11566 16507
rect 11882 16504 11888 16516
rect 11554 16476 11888 16504
rect 11554 16473 11566 16476
rect 11508 16467 11566 16473
rect 11882 16464 11888 16476
rect 11940 16464 11946 16516
rect 14277 16507 14335 16513
rect 14277 16473 14289 16507
rect 14323 16504 14335 16507
rect 14366 16504 14372 16516
rect 14323 16476 14372 16504
rect 14323 16473 14335 16476
rect 14277 16467 14335 16473
rect 14366 16464 14372 16476
rect 14424 16464 14430 16516
rect 7374 16436 7380 16448
rect 5828 16408 7380 16436
rect 7374 16396 7380 16408
rect 7432 16436 7438 16448
rect 8389 16439 8447 16445
rect 8389 16436 8401 16439
rect 7432 16408 8401 16436
rect 7432 16396 7438 16408
rect 8389 16405 8401 16408
rect 8435 16405 8447 16439
rect 8389 16399 8447 16405
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 12621 16439 12679 16445
rect 12621 16436 12633 16439
rect 12492 16408 12633 16436
rect 12492 16396 12498 16408
rect 12621 16405 12633 16408
rect 12667 16405 12679 16439
rect 14826 16436 14832 16448
rect 14787 16408 14832 16436
rect 12621 16399 12679 16405
rect 14826 16396 14832 16408
rect 14884 16396 14890 16448
rect 16025 16439 16083 16445
rect 16025 16405 16037 16439
rect 16071 16436 16083 16439
rect 16298 16436 16304 16448
rect 16071 16408 16304 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 1104 16346 18860 16368
rect 1104 16294 6880 16346
rect 6932 16294 6944 16346
rect 6996 16294 7008 16346
rect 7060 16294 7072 16346
rect 7124 16294 7136 16346
rect 7188 16294 12811 16346
rect 12863 16294 12875 16346
rect 12927 16294 12939 16346
rect 12991 16294 13003 16346
rect 13055 16294 13067 16346
rect 13119 16294 18860 16346
rect 1104 16272 18860 16294
rect 2958 16192 2964 16244
rect 3016 16232 3022 16244
rect 3697 16235 3755 16241
rect 3697 16232 3709 16235
rect 3016 16204 3709 16232
rect 3016 16192 3022 16204
rect 3697 16201 3709 16204
rect 3743 16201 3755 16235
rect 6730 16232 6736 16244
rect 6691 16204 6736 16232
rect 3697 16195 3755 16201
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 10962 16232 10968 16244
rect 8628 16204 9996 16232
rect 10923 16204 10968 16232
rect 8628 16192 8634 16204
rect 2593 16167 2651 16173
rect 2593 16133 2605 16167
rect 2639 16133 2651 16167
rect 2593 16127 2651 16133
rect 2608 16096 2636 16127
rect 2774 16124 2780 16176
rect 2832 16173 2838 16176
rect 2832 16167 2851 16173
rect 2839 16133 2851 16167
rect 2832 16127 2851 16133
rect 2832 16124 2838 16127
rect 6178 16124 6184 16176
rect 6236 16164 6242 16176
rect 6365 16167 6423 16173
rect 6365 16164 6377 16167
rect 6236 16136 6377 16164
rect 6236 16124 6242 16136
rect 6365 16133 6377 16136
rect 6411 16133 6423 16167
rect 6365 16127 6423 16133
rect 6581 16167 6639 16173
rect 6581 16133 6593 16167
rect 6627 16164 6639 16167
rect 7282 16164 7288 16176
rect 6627 16136 7288 16164
rect 6627 16133 6639 16136
rect 6581 16127 6639 16133
rect 3234 16096 3240 16108
rect 2608 16068 3240 16096
rect 3234 16056 3240 16068
rect 3292 16096 3298 16108
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 3292 16068 3985 16096
rect 3292 16056 3298 16068
rect 3973 16065 3985 16068
rect 4019 16096 4031 16099
rect 4154 16096 4160 16108
rect 4019 16068 4160 16096
rect 4019 16065 4031 16068
rect 3973 16059 4031 16065
rect 4154 16056 4160 16068
rect 4212 16096 4218 16108
rect 5442 16096 5448 16108
rect 4212 16068 5448 16096
rect 4212 16056 4218 16068
rect 5442 16056 5448 16068
rect 5500 16096 5506 16108
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 5500 16068 5549 16096
rect 5500 16056 5506 16068
rect 5537 16065 5549 16068
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5776 16068 5825 16096
rect 5776 16056 5782 16068
rect 5813 16065 5825 16068
rect 5859 16065 5871 16099
rect 6380 16096 6408 16127
rect 7282 16124 7288 16136
rect 7340 16124 7346 16176
rect 7834 16124 7840 16176
rect 7892 16164 7898 16176
rect 8110 16164 8116 16176
rect 7892 16136 8116 16164
rect 7892 16124 7898 16136
rect 8110 16124 8116 16136
rect 8168 16164 8174 16176
rect 8168 16136 8708 16164
rect 8168 16124 8174 16136
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 6380 16068 7757 16096
rect 5813 16059 5871 16065
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 8018 16096 8024 16108
rect 7979 16068 8024 16096
rect 7745 16059 7803 16065
rect 8018 16056 8024 16068
rect 8076 16096 8082 16108
rect 8680 16105 8708 16136
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 9968 16173 9996 16204
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 11977 16235 12035 16241
rect 11977 16201 11989 16235
rect 12023 16232 12035 16235
rect 12066 16232 12072 16244
rect 12023 16204 12072 16232
rect 12023 16201 12035 16204
rect 11977 16195 12035 16201
rect 12066 16192 12072 16204
rect 12124 16192 12130 16244
rect 17310 16232 17316 16244
rect 17271 16204 17316 16232
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 9861 16167 9919 16173
rect 9861 16164 9873 16167
rect 9732 16136 9873 16164
rect 9732 16124 9738 16136
rect 9861 16133 9873 16136
rect 9907 16133 9919 16167
rect 9861 16127 9919 16133
rect 9953 16167 10011 16173
rect 9953 16133 9965 16167
rect 9999 16133 10011 16167
rect 9953 16127 10011 16133
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 10284 16136 10824 16164
rect 10284 16124 10290 16136
rect 8481 16099 8539 16105
rect 8481 16096 8493 16099
rect 8076 16068 8493 16096
rect 8076 16056 8082 16068
rect 8481 16065 8493 16068
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16065 8723 16099
rect 8665 16059 8723 16065
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16065 8999 16099
rect 9766 16096 9772 16108
rect 9727 16068 9772 16096
rect 8941 16059 8999 16065
rect 3050 15988 3056 16040
rect 3108 16028 3114 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3108 16000 3433 16028
rect 3108 15988 3114 16000
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 3694 15988 3700 16040
rect 3752 16028 3758 16040
rect 4065 16031 4123 16037
rect 4065 16028 4077 16031
rect 3752 16000 4077 16028
rect 3752 15988 3758 16000
rect 4065 15997 4077 16000
rect 4111 15997 4123 16031
rect 8956 16028 8984 16059
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 10134 16096 10140 16108
rect 10095 16068 10140 16096
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 10686 16096 10692 16108
rect 10647 16068 10692 16096
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 10796 16105 10824 16136
rect 12342 16124 12348 16176
rect 12400 16164 12406 16176
rect 12400 16136 13400 16164
rect 12400 16124 12406 16136
rect 13372 16105 13400 16136
rect 10781 16099 10839 16105
rect 10781 16065 10793 16099
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 13101 16099 13159 16105
rect 13101 16065 13113 16099
rect 13147 16096 13159 16099
rect 13357 16099 13415 16105
rect 13147 16068 13308 16096
rect 13147 16065 13159 16068
rect 13101 16059 13159 16065
rect 10410 16028 10416 16040
rect 8956 16000 10416 16028
rect 4065 15991 4123 15997
rect 10410 15988 10416 16000
rect 10468 15988 10474 16040
rect 13280 16028 13308 16068
rect 13357 16065 13369 16099
rect 13403 16065 13415 16099
rect 17494 16096 17500 16108
rect 17455 16068 17500 16096
rect 13357 16059 13415 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 14826 16028 14832 16040
rect 13280 16000 14832 16028
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 3068 15960 3096 15988
rect 2792 15932 3096 15960
rect 2792 15901 2820 15932
rect 3326 15920 3332 15972
rect 3384 15960 3390 15972
rect 6086 15960 6092 15972
rect 3384 15932 6092 15960
rect 3384 15920 3390 15932
rect 6086 15920 6092 15932
rect 6144 15920 6150 15972
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15861 2835 15895
rect 2777 15855 2835 15861
rect 2961 15895 3019 15901
rect 2961 15861 2973 15895
rect 3007 15892 3019 15895
rect 3418 15892 3424 15904
rect 3007 15864 3424 15892
rect 3007 15861 3019 15864
rect 2961 15855 3019 15861
rect 3418 15852 3424 15864
rect 3476 15852 3482 15904
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 8444 15864 9137 15892
rect 8444 15852 8450 15864
rect 9125 15861 9137 15864
rect 9171 15861 9183 15895
rect 9582 15892 9588 15904
rect 9543 15864 9588 15892
rect 9125 15855 9183 15861
rect 9582 15852 9588 15864
rect 9640 15852 9646 15904
rect 1104 15802 18860 15824
rect 1104 15750 3915 15802
rect 3967 15750 3979 15802
rect 4031 15750 4043 15802
rect 4095 15750 4107 15802
rect 4159 15750 4171 15802
rect 4223 15750 9846 15802
rect 9898 15750 9910 15802
rect 9962 15750 9974 15802
rect 10026 15750 10038 15802
rect 10090 15750 10102 15802
rect 10154 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 15904 15802
rect 15956 15750 15968 15802
rect 16020 15750 16032 15802
rect 16084 15750 18860 15802
rect 1104 15728 18860 15750
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 6089 15691 6147 15697
rect 6089 15657 6101 15691
rect 6135 15688 6147 15691
rect 6454 15688 6460 15700
rect 6135 15660 6460 15688
rect 6135 15657 6147 15660
rect 6089 15651 6147 15657
rect 6454 15648 6460 15660
rect 6512 15648 6518 15700
rect 7745 15691 7803 15697
rect 7745 15657 7757 15691
rect 7791 15688 7803 15691
rect 8202 15688 8208 15700
rect 7791 15660 8208 15688
rect 7791 15657 7803 15660
rect 7745 15651 7803 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 11517 15691 11575 15697
rect 11517 15688 11529 15691
rect 11020 15660 11529 15688
rect 11020 15648 11026 15660
rect 11517 15657 11529 15660
rect 11563 15657 11575 15691
rect 11517 15651 11575 15657
rect 3237 15623 3295 15629
rect 3237 15589 3249 15623
rect 3283 15620 3295 15623
rect 3326 15620 3332 15632
rect 3283 15592 3332 15620
rect 3283 15589 3295 15592
rect 3237 15583 3295 15589
rect 3326 15580 3332 15592
rect 3384 15580 3390 15632
rect 7650 15620 7656 15632
rect 5828 15592 7656 15620
rect 3786 15512 3792 15564
rect 3844 15552 3850 15564
rect 3881 15555 3939 15561
rect 3881 15552 3893 15555
rect 3844 15524 3893 15552
rect 3844 15512 3850 15524
rect 3881 15521 3893 15524
rect 3927 15521 3939 15555
rect 3881 15515 3939 15521
rect 2774 15444 2780 15496
rect 2832 15484 2838 15496
rect 2961 15487 3019 15493
rect 2961 15484 2973 15487
rect 2832 15456 2973 15484
rect 2832 15444 2838 15456
rect 2961 15453 2973 15456
rect 3007 15484 3019 15487
rect 3694 15484 3700 15496
rect 3007 15456 3700 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 5828 15493 5856 15592
rect 7650 15580 7656 15592
rect 7708 15580 7714 15632
rect 8294 15620 8300 15632
rect 7944 15592 8300 15620
rect 6546 15552 6552 15564
rect 6507 15524 6552 15552
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15552 7251 15555
rect 7282 15552 7288 15564
rect 7239 15524 7288 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 5905 15487 5963 15493
rect 5905 15453 5917 15487
rect 5951 15484 5963 15487
rect 6178 15484 6184 15496
rect 5951 15456 6184 15484
rect 5951 15453 5963 15456
rect 5905 15447 5963 15453
rect 6178 15444 6184 15456
rect 6236 15484 6242 15496
rect 7944 15493 7972 15592
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 8018 15512 8024 15564
rect 8076 15512 8082 15564
rect 10965 15555 11023 15561
rect 10965 15521 10977 15555
rect 11011 15552 11023 15555
rect 11238 15552 11244 15564
rect 11011 15524 11244 15552
rect 11011 15521 11023 15524
rect 10965 15515 11023 15521
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 11701 15555 11759 15561
rect 11701 15552 11713 15555
rect 11388 15524 11713 15552
rect 11388 15512 11394 15524
rect 11701 15521 11713 15524
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 7101 15487 7159 15493
rect 7101 15484 7113 15487
rect 6236 15456 7113 15484
rect 6236 15444 6242 15456
rect 7101 15453 7113 15456
rect 7147 15453 7159 15487
rect 7101 15447 7159 15453
rect 7924 15487 7982 15493
rect 7924 15453 7936 15487
rect 7970 15453 7982 15487
rect 8036 15484 8064 15512
rect 8241 15487 8299 15493
rect 8241 15484 8253 15487
rect 8036 15456 8253 15484
rect 7924 15447 7982 15453
rect 8241 15453 8253 15456
rect 8287 15453 8299 15487
rect 8241 15447 8299 15453
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 11425 15487 11483 15493
rect 8444 15456 8489 15484
rect 8444 15444 8450 15456
rect 11425 15453 11437 15487
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 12345 15487 12403 15493
rect 12345 15453 12357 15487
rect 12391 15484 12403 15487
rect 12526 15484 12532 15496
rect 12391 15456 12532 15484
rect 12391 15453 12403 15456
rect 12345 15447 12403 15453
rect 3234 15416 3240 15428
rect 3195 15388 3240 15416
rect 3234 15376 3240 15388
rect 3292 15376 3298 15428
rect 4148 15419 4206 15425
rect 4148 15385 4160 15419
rect 4194 15416 4206 15419
rect 4246 15416 4252 15428
rect 4194 15388 4252 15416
rect 4194 15385 4206 15388
rect 4148 15379 4206 15385
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 6086 15416 6092 15428
rect 6047 15388 6092 15416
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 7374 15376 7380 15428
rect 7432 15416 7438 15428
rect 8021 15419 8079 15425
rect 8021 15416 8033 15419
rect 7432 15388 8033 15416
rect 7432 15376 7438 15388
rect 8021 15385 8033 15388
rect 8067 15385 8079 15419
rect 8021 15379 8079 15385
rect 8110 15376 8116 15428
rect 8168 15416 8174 15428
rect 10720 15419 10778 15425
rect 8168 15388 8213 15416
rect 8168 15376 8174 15388
rect 10720 15385 10732 15419
rect 10766 15416 10778 15419
rect 10870 15416 10876 15428
rect 10766 15388 10876 15416
rect 10766 15385 10778 15388
rect 10720 15379 10778 15385
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 3050 15348 3056 15360
rect 3011 15320 3056 15348
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 6730 15308 6736 15360
rect 6788 15348 6794 15360
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 6788 15320 6837 15348
rect 6788 15308 6794 15320
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 9585 15351 9643 15357
rect 9585 15317 9597 15351
rect 9631 15348 9643 15351
rect 10318 15348 10324 15360
rect 9631 15320 10324 15348
rect 9631 15317 9643 15320
rect 9585 15311 9643 15317
rect 10318 15308 10324 15320
rect 10376 15348 10382 15360
rect 11440 15348 11468 15447
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 12066 15376 12072 15428
rect 12124 15416 12130 15428
rect 14185 15419 14243 15425
rect 14185 15416 14197 15419
rect 12124 15388 14197 15416
rect 12124 15376 12130 15388
rect 14185 15385 14197 15388
rect 14231 15385 14243 15419
rect 14366 15416 14372 15428
rect 14327 15388 14372 15416
rect 14185 15379 14243 15385
rect 14366 15376 14372 15388
rect 14424 15376 14430 15428
rect 11698 15348 11704 15360
rect 10376 15320 11468 15348
rect 11659 15320 11704 15348
rect 10376 15308 10382 15320
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 11882 15308 11888 15360
rect 11940 15348 11946 15360
rect 12161 15351 12219 15357
rect 12161 15348 12173 15351
rect 11940 15320 12173 15348
rect 11940 15308 11946 15320
rect 12161 15317 12173 15320
rect 12207 15317 12219 15351
rect 12161 15311 12219 15317
rect 1104 15258 18860 15280
rect 1104 15206 6880 15258
rect 6932 15206 6944 15258
rect 6996 15206 7008 15258
rect 7060 15206 7072 15258
rect 7124 15206 7136 15258
rect 7188 15206 12811 15258
rect 12863 15206 12875 15258
rect 12927 15206 12939 15258
rect 12991 15206 13003 15258
rect 13055 15206 13067 15258
rect 13119 15206 18860 15258
rect 1104 15184 18860 15206
rect 3602 15144 3608 15156
rect 3563 15116 3608 15144
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 3694 15104 3700 15156
rect 3752 15144 3758 15156
rect 4065 15147 4123 15153
rect 4065 15144 4077 15147
rect 3752 15116 4077 15144
rect 3752 15104 3758 15116
rect 4065 15113 4077 15116
rect 4111 15113 4123 15147
rect 4065 15107 4123 15113
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 7561 15147 7619 15153
rect 7561 15144 7573 15147
rect 6604 15116 7573 15144
rect 6604 15104 6610 15116
rect 7561 15113 7573 15116
rect 7607 15113 7619 15147
rect 7561 15107 7619 15113
rect 10121 15147 10179 15153
rect 10121 15113 10133 15147
rect 10167 15144 10179 15147
rect 10226 15144 10232 15156
rect 10167 15116 10232 15144
rect 10167 15113 10179 15116
rect 10121 15107 10179 15113
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 10870 15144 10876 15156
rect 10831 15116 10876 15144
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 4246 15076 4252 15088
rect 4159 15048 4252 15076
rect 4246 15036 4252 15048
rect 4304 15076 4310 15088
rect 5258 15076 5264 15088
rect 4304 15048 5264 15076
rect 4304 15036 4310 15048
rect 5258 15036 5264 15048
rect 5316 15036 5322 15088
rect 8386 15036 8392 15088
rect 8444 15076 8450 15088
rect 9674 15076 9680 15088
rect 8444 15048 9680 15076
rect 8444 15036 8450 15048
rect 3326 15008 3332 15020
rect 3287 14980 3332 15008
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 3418 14968 3424 15020
rect 3476 15008 3482 15020
rect 4430 15008 4436 15020
rect 3476 14980 3521 15008
rect 4391 14980 4436 15008
rect 3476 14968 3482 14980
rect 4430 14968 4436 14980
rect 4488 14968 4494 15020
rect 6914 15008 6920 15020
rect 6875 14980 6920 15008
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 7432 14980 7573 15008
rect 7432 14968 7438 14980
rect 7561 14977 7573 14980
rect 7607 14977 7619 15011
rect 7742 15008 7748 15020
rect 7703 14980 7748 15008
rect 7561 14971 7619 14977
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 8570 15008 8576 15020
rect 8531 14980 8576 15008
rect 8570 14968 8576 14980
rect 8628 14968 8634 15020
rect 8864 15017 8892 15048
rect 9674 15036 9680 15048
rect 9732 15036 9738 15088
rect 10318 15076 10324 15088
rect 10279 15048 10324 15076
rect 10318 15036 10324 15048
rect 10376 15036 10382 15088
rect 11974 15076 11980 15088
rect 11935 15048 11980 15076
rect 11974 15036 11980 15048
rect 12032 15036 12038 15088
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 15008 8999 15011
rect 9766 15008 9772 15020
rect 8987 14980 9772 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 10226 14968 10232 15020
rect 10284 15008 10290 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10284 14980 10793 15008
rect 10284 14968 10290 14980
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 15008 11023 15011
rect 11698 15008 11704 15020
rect 11011 14980 11704 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 17681 15011 17739 15017
rect 17681 14977 17693 15011
rect 17727 15008 17739 15011
rect 17954 15008 17960 15020
rect 17727 14980 17960 15008
rect 17727 14977 17739 14980
rect 17681 14971 17739 14977
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 3510 14900 3516 14952
rect 3568 14940 3574 14952
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3568 14912 3617 14940
rect 3568 14900 3574 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 8665 14943 8723 14949
rect 8665 14909 8677 14943
rect 8711 14940 8723 14943
rect 9214 14940 9220 14952
rect 8711 14912 9220 14940
rect 8711 14909 8723 14912
rect 8665 14903 8723 14909
rect 9214 14900 9220 14912
rect 9272 14940 9278 14952
rect 9490 14940 9496 14952
rect 9272 14912 9496 14940
rect 9272 14900 9278 14912
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 17862 14940 17868 14952
rect 17823 14912 17868 14940
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 7101 14875 7159 14881
rect 7101 14841 7113 14875
rect 7147 14872 7159 14875
rect 7650 14872 7656 14884
rect 7147 14844 7656 14872
rect 7147 14841 7159 14844
rect 7101 14835 7159 14841
rect 7650 14832 7656 14844
rect 7708 14832 7714 14884
rect 9953 14875 10011 14881
rect 9953 14841 9965 14875
rect 9999 14872 10011 14875
rect 10226 14872 10232 14884
rect 9999 14844 10232 14872
rect 9999 14841 10011 14844
rect 9953 14835 10011 14841
rect 10226 14832 10232 14844
rect 10284 14832 10290 14884
rect 9122 14804 9128 14816
rect 9083 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 10137 14807 10195 14813
rect 10137 14773 10149 14807
rect 10183 14804 10195 14807
rect 10686 14804 10692 14816
rect 10183 14776 10692 14804
rect 10183 14773 10195 14776
rect 10137 14767 10195 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 12066 14804 12072 14816
rect 12027 14776 12072 14804
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 1104 14714 18860 14736
rect 1104 14662 3915 14714
rect 3967 14662 3979 14714
rect 4031 14662 4043 14714
rect 4095 14662 4107 14714
rect 4159 14662 4171 14714
rect 4223 14662 9846 14714
rect 9898 14662 9910 14714
rect 9962 14662 9974 14714
rect 10026 14662 10038 14714
rect 10090 14662 10102 14714
rect 10154 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 15904 14714
rect 15956 14662 15968 14714
rect 16020 14662 16032 14714
rect 16084 14662 18860 14714
rect 1104 14640 18860 14662
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3108 14572 4077 14600
rect 3108 14560 3114 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 8996 14572 9321 14600
rect 8996 14560 9002 14572
rect 9309 14569 9321 14572
rect 9355 14569 9367 14603
rect 17954 14600 17960 14612
rect 17915 14572 17960 14600
rect 9309 14563 9367 14569
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 6914 14492 6920 14544
rect 6972 14532 6978 14544
rect 7834 14532 7840 14544
rect 6972 14504 7840 14532
rect 6972 14492 6978 14504
rect 7834 14492 7840 14504
rect 7892 14532 7898 14544
rect 13538 14532 13544 14544
rect 7892 14504 13544 14532
rect 7892 14492 7898 14504
rect 13538 14492 13544 14504
rect 13596 14492 13602 14544
rect 9401 14467 9459 14473
rect 9401 14433 9413 14467
rect 9447 14464 9459 14467
rect 9582 14464 9588 14476
rect 9447 14436 9588 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 11514 14464 11520 14476
rect 9692 14436 11520 14464
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4246 14396 4252 14408
rect 4203 14368 4252 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 3988 14328 4016 14359
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 9122 14396 9128 14408
rect 9083 14368 9128 14396
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 4430 14328 4436 14340
rect 3988 14300 4436 14328
rect 4430 14288 4436 14300
rect 4488 14328 4494 14340
rect 9692 14328 9720 14436
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 10686 14396 10692 14408
rect 10643 14368 10692 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15620 14368 15761 14396
rect 15620 14356 15626 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 18138 14396 18144 14408
rect 18099 14368 18144 14396
rect 15749 14359 15807 14365
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 9858 14328 9864 14340
rect 4488 14300 9720 14328
rect 9819 14300 9864 14328
rect 4488 14288 4494 14300
rect 9858 14288 9864 14300
rect 9916 14288 9922 14340
rect 10045 14331 10103 14337
rect 10045 14297 10057 14331
rect 10091 14328 10103 14331
rect 12066 14328 12072 14340
rect 10091 14300 12072 14328
rect 10091 14297 10103 14300
rect 10045 14291 10103 14297
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 8938 14260 8944 14272
rect 8899 14232 8944 14260
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 10689 14263 10747 14269
rect 10689 14260 10701 14263
rect 9732 14232 10701 14260
rect 9732 14220 9738 14232
rect 10689 14229 10701 14232
rect 10735 14229 10747 14263
rect 10689 14223 10747 14229
rect 15010 14220 15016 14272
rect 15068 14260 15074 14272
rect 15565 14263 15623 14269
rect 15565 14260 15577 14263
rect 15068 14232 15577 14260
rect 15068 14220 15074 14232
rect 15565 14229 15577 14232
rect 15611 14229 15623 14263
rect 15565 14223 15623 14229
rect 1104 14170 18860 14192
rect 1104 14118 6880 14170
rect 6932 14118 6944 14170
rect 6996 14118 7008 14170
rect 7060 14118 7072 14170
rect 7124 14118 7136 14170
rect 7188 14118 12811 14170
rect 12863 14118 12875 14170
rect 12927 14118 12939 14170
rect 12991 14118 13003 14170
rect 13055 14118 13067 14170
rect 13119 14118 18860 14170
rect 1104 14096 18860 14118
rect 15562 14056 15568 14068
rect 15523 14028 15568 14056
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 9585 13991 9643 13997
rect 9585 13988 9597 13991
rect 9364 13960 9597 13988
rect 9364 13948 9370 13960
rect 9585 13957 9597 13960
rect 9631 13957 9643 13991
rect 9585 13951 9643 13957
rect 9769 13991 9827 13997
rect 9769 13957 9781 13991
rect 9815 13988 9827 13991
rect 9858 13988 9864 14000
rect 9815 13960 9864 13988
rect 9815 13957 9827 13960
rect 9769 13951 9827 13957
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 14366 13948 14372 14000
rect 14424 13988 14430 14000
rect 14553 13991 14611 13997
rect 14553 13988 14565 13991
rect 14424 13960 14565 13988
rect 14424 13948 14430 13960
rect 14553 13957 14565 13960
rect 14599 13957 14611 13991
rect 14553 13951 14611 13957
rect 13814 13920 13820 13932
rect 13775 13892 13820 13920
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 15749 13923 15807 13929
rect 15749 13889 15761 13923
rect 15795 13920 15807 13923
rect 16390 13920 16396 13932
rect 15795 13892 16396 13920
rect 15795 13889 15807 13892
rect 15749 13883 15807 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 13633 13855 13691 13861
rect 13633 13852 13645 13855
rect 13412 13824 13645 13852
rect 13412 13812 13418 13824
rect 13633 13821 13645 13824
rect 13679 13821 13691 13855
rect 13633 13815 13691 13821
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14458 13852 14464 13864
rect 14047 13824 14464 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 15654 13812 15660 13864
rect 15712 13852 15718 13864
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 15712 13824 15945 13852
rect 15712 13812 15718 13824
rect 15933 13821 15945 13824
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 14734 13784 14740 13796
rect 14695 13756 14740 13784
rect 14734 13744 14740 13756
rect 14792 13744 14798 13796
rect 1104 13626 18860 13648
rect 1104 13574 3915 13626
rect 3967 13574 3979 13626
rect 4031 13574 4043 13626
rect 4095 13574 4107 13626
rect 4159 13574 4171 13626
rect 4223 13574 9846 13626
rect 9898 13574 9910 13626
rect 9962 13574 9974 13626
rect 10026 13574 10038 13626
rect 10090 13574 10102 13626
rect 10154 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 15904 13626
rect 15956 13574 15968 13626
rect 16020 13574 16032 13626
rect 16084 13574 18860 13626
rect 1104 13552 18860 13574
rect 15933 13515 15991 13521
rect 15933 13481 15945 13515
rect 15979 13512 15991 13515
rect 16114 13512 16120 13524
rect 15979 13484 16120 13512
rect 15979 13481 15991 13484
rect 15933 13475 15991 13481
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 16298 13472 16304 13524
rect 16356 13512 16362 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 16356 13484 16957 13512
rect 16356 13472 16362 13484
rect 16945 13481 16957 13484
rect 16991 13481 17003 13515
rect 17402 13512 17408 13524
rect 17363 13484 17408 13512
rect 16945 13475 17003 13481
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 16206 13336 16212 13388
rect 16264 13376 16270 13388
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 16264 13348 17049 13376
rect 16264 13336 16270 13348
rect 17037 13345 17049 13348
rect 17083 13345 17095 13379
rect 17037 13339 17095 13345
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13538 13308 13544 13320
rect 13403 13280 13544 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 13280 13240 13308 13271
rect 13538 13268 13544 13280
rect 13596 13308 13602 13320
rect 13814 13308 13820 13320
rect 13596 13280 13820 13308
rect 13596 13268 13602 13280
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 14792 13280 15485 13308
rect 14792 13268 14798 13280
rect 15473 13277 15485 13280
rect 15519 13277 15531 13311
rect 16298 13308 16304 13320
rect 16259 13280 16304 13308
rect 15473 13271 15531 13277
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13308 16543 13311
rect 16666 13308 16672 13320
rect 16531 13280 16672 13308
rect 16531 13277 16543 13280
rect 16485 13271 16543 13277
rect 16666 13268 16672 13280
rect 16724 13308 16730 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 16724 13280 17233 13308
rect 16724 13268 16730 13280
rect 17221 13277 17233 13280
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 13446 13240 13452 13252
rect 13280 13212 13452 13240
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 14642 13200 14648 13252
rect 14700 13240 14706 13252
rect 15206 13243 15264 13249
rect 15206 13240 15218 13243
rect 14700 13212 15218 13240
rect 14700 13200 14706 13212
rect 15206 13209 15218 13212
rect 15252 13209 15264 13243
rect 15206 13203 15264 13209
rect 15654 13200 15660 13252
rect 15712 13240 15718 13252
rect 16117 13243 16175 13249
rect 16117 13240 16129 13243
rect 15712 13212 16129 13240
rect 15712 13200 15718 13212
rect 16117 13209 16129 13212
rect 16163 13240 16175 13243
rect 16945 13243 17003 13249
rect 16945 13240 16957 13243
rect 16163 13212 16957 13240
rect 16163 13209 16175 13212
rect 16117 13203 16175 13209
rect 16945 13209 16957 13212
rect 16991 13209 17003 13243
rect 16945 13203 17003 13209
rect 13541 13175 13599 13181
rect 13541 13141 13553 13175
rect 13587 13172 13599 13175
rect 13814 13172 13820 13184
rect 13587 13144 13820 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 14090 13172 14096 13184
rect 14051 13144 14096 13172
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 16206 13172 16212 13184
rect 16167 13144 16212 13172
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 1104 13082 18860 13104
rect 1104 13030 6880 13082
rect 6932 13030 6944 13082
rect 6996 13030 7008 13082
rect 7060 13030 7072 13082
rect 7124 13030 7136 13082
rect 7188 13030 12811 13082
rect 12863 13030 12875 13082
rect 12927 13030 12939 13082
rect 12991 13030 13003 13082
rect 13055 13030 13067 13082
rect 13119 13030 18860 13082
rect 1104 13008 18860 13030
rect 12989 12971 13047 12977
rect 12989 12937 13001 12971
rect 13035 12968 13047 12971
rect 13262 12968 13268 12980
rect 13035 12940 13268 12968
rect 13035 12937 13047 12940
rect 12989 12931 13047 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 8570 12900 8576 12912
rect 8531 12872 8576 12900
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 9585 12903 9643 12909
rect 9585 12869 9597 12903
rect 9631 12900 9643 12903
rect 9766 12900 9772 12912
rect 9631 12872 9772 12900
rect 9631 12869 9643 12872
rect 9585 12863 9643 12869
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 16117 12903 16175 12909
rect 16117 12869 16129 12903
rect 16163 12900 16175 12903
rect 16163 12872 17724 12900
rect 16163 12869 16175 12872
rect 16117 12863 16175 12869
rect 10318 12832 10324 12844
rect 10279 12804 10324 12832
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 11876 12835 11934 12841
rect 11876 12801 11888 12835
rect 11922 12832 11934 12835
rect 13722 12832 13728 12844
rect 11922 12804 13728 12832
rect 11922 12801 11934 12804
rect 11876 12795 11934 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14562 12835 14620 12841
rect 14562 12832 14574 12835
rect 14332 12804 14574 12832
rect 14332 12792 14338 12804
rect 14562 12801 14574 12804
rect 14608 12801 14620 12835
rect 14562 12795 14620 12801
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 14792 12804 14841 12832
rect 14792 12792 14798 12804
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16390 12832 16396 12844
rect 15979 12804 16396 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16390 12792 16396 12804
rect 16448 12832 16454 12844
rect 17696 12841 17724 12872
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16448 12804 16865 12832
rect 16448 12792 16454 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12801 17739 12835
rect 17681 12795 17739 12801
rect 11606 12764 11612 12776
rect 11567 12736 11612 12764
rect 11606 12724 11612 12736
rect 11664 12724 11670 12776
rect 15749 12767 15807 12773
rect 15749 12733 15761 12767
rect 15795 12764 15807 12767
rect 16298 12764 16304 12776
rect 15795 12736 16304 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16666 12724 16672 12776
rect 16724 12764 16730 12776
rect 16724 12736 16769 12764
rect 16724 12724 16730 12736
rect 8662 12628 8668 12640
rect 8623 12600 8668 12628
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 9493 12631 9551 12637
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 9582 12628 9588 12640
rect 9539 12600 9588 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10229 12631 10287 12637
rect 10229 12628 10241 12631
rect 9824 12600 10241 12628
rect 9824 12588 9830 12600
rect 10229 12597 10241 12600
rect 10275 12597 10287 12631
rect 10229 12591 10287 12597
rect 13354 12588 13360 12640
rect 13412 12628 13418 12640
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 13412 12600 13461 12628
rect 13412 12588 13418 12600
rect 13449 12597 13461 12600
rect 13495 12597 13507 12631
rect 13449 12591 13507 12597
rect 17037 12631 17095 12637
rect 17037 12597 17049 12631
rect 17083 12628 17095 12631
rect 17402 12628 17408 12640
rect 17083 12600 17408 12628
rect 17083 12597 17095 12600
rect 17037 12591 17095 12597
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 17494 12588 17500 12640
rect 17552 12628 17558 12640
rect 17552 12600 17597 12628
rect 17552 12588 17558 12600
rect 1104 12538 18860 12560
rect 1104 12486 3915 12538
rect 3967 12486 3979 12538
rect 4031 12486 4043 12538
rect 4095 12486 4107 12538
rect 4159 12486 4171 12538
rect 4223 12486 9846 12538
rect 9898 12486 9910 12538
rect 9962 12486 9974 12538
rect 10026 12486 10038 12538
rect 10090 12486 10102 12538
rect 10154 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 15904 12538
rect 15956 12486 15968 12538
rect 16020 12486 16032 12538
rect 16084 12486 18860 12538
rect 1104 12464 18860 12486
rect 8389 12427 8447 12433
rect 8389 12393 8401 12427
rect 8435 12424 8447 12427
rect 8570 12424 8576 12436
rect 8435 12396 8576 12424
rect 8435 12393 8447 12396
rect 8389 12387 8447 12393
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 12710 12424 12716 12436
rect 12391 12396 12716 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13780 12396 14105 12424
rect 13780 12384 13786 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14240 12396 14504 12424
rect 14240 12384 14246 12396
rect 9030 12316 9036 12368
rect 9088 12356 9094 12368
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 9088 12328 10057 12356
rect 9088 12316 9094 12328
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 10045 12319 10103 12325
rect 13541 12359 13599 12365
rect 13541 12325 13553 12359
rect 13587 12356 13599 12359
rect 13587 12328 14412 12356
rect 13587 12325 13599 12328
rect 13541 12319 13599 12325
rect 9582 12288 9588 12300
rect 8864 12260 9588 12288
rect 8864 12232 8892 12260
rect 9582 12248 9588 12260
rect 9640 12288 9646 12300
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 9640 12260 10977 12288
rect 9640 12248 9646 12260
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 3844 12192 7021 12220
rect 3844 12180 3850 12192
rect 7009 12189 7021 12192
rect 7055 12220 7067 12223
rect 8846 12220 8852 12232
rect 7055 12192 8852 12220
rect 7055 12189 7067 12192
rect 7009 12183 7067 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 9089 12223 9147 12229
rect 8996 12192 9041 12220
rect 8996 12180 9002 12192
rect 9089 12189 9101 12223
rect 9135 12220 9147 12223
rect 9135 12189 9168 12220
rect 9089 12183 9168 12189
rect 7282 12161 7288 12164
rect 7276 12115 7288 12161
rect 7340 12152 7346 12164
rect 7340 12124 7376 12152
rect 7282 12112 7288 12115
rect 7340 12112 7346 12124
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 9140 12152 9168 12183
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9447 12223 9505 12229
rect 9272 12192 9317 12220
rect 9272 12180 9278 12192
rect 9447 12189 9459 12223
rect 9493 12220 9505 12223
rect 9766 12220 9772 12232
rect 9493 12192 9772 12220
rect 9493 12189 9505 12192
rect 9447 12183 9505 12189
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 10192 12192 10333 12220
rect 10192 12180 10198 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10980 12220 11008 12251
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 14182 12288 14188 12300
rect 12216 12260 14188 12288
rect 12216 12248 12222 12260
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 11606 12220 11612 12232
rect 10980 12192 11612 12220
rect 10321 12183 10379 12189
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12220 13323 12223
rect 14090 12220 14096 12232
rect 13311 12192 14096 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14384 12229 14412 12328
rect 14476 12229 14504 12396
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 16724 12396 16773 12424
rect 16724 12384 16730 12396
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 16761 12387 16819 12393
rect 14734 12316 14740 12368
rect 14792 12316 14798 12368
rect 14752 12288 14780 12316
rect 15381 12291 15439 12297
rect 15381 12288 15393 12291
rect 14752 12260 15393 12288
rect 15381 12257 15393 12260
rect 15427 12257 15439 12291
rect 15381 12251 15439 12257
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 14200 12192 14289 12220
rect 9306 12152 9312 12164
rect 8720 12124 9168 12152
rect 9267 12124 9312 12152
rect 8720 12112 8726 12124
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 10045 12155 10103 12161
rect 10045 12121 10057 12155
rect 10091 12152 10103 12155
rect 10502 12152 10508 12164
rect 10091 12124 10508 12152
rect 10091 12121 10103 12124
rect 10045 12115 10103 12121
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 11232 12155 11290 12161
rect 11232 12121 11244 12155
rect 11278 12152 11290 12155
rect 11790 12152 11796 12164
rect 11278 12124 11796 12152
rect 11278 12121 11290 12124
rect 11232 12115 11290 12121
rect 11790 12112 11796 12124
rect 11848 12112 11854 12164
rect 12989 12155 13047 12161
rect 12989 12121 13001 12155
rect 13035 12152 13047 12155
rect 13446 12152 13452 12164
rect 13035 12124 13452 12152
rect 13035 12121 13047 12124
rect 12989 12115 13047 12121
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 9585 12087 9643 12093
rect 9585 12053 9597 12087
rect 9631 12084 9643 12087
rect 9674 12084 9680 12096
rect 9631 12056 9680 12084
rect 9631 12053 9643 12056
rect 9585 12047 9643 12053
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 10229 12087 10287 12093
rect 10229 12053 10241 12087
rect 10275 12084 10287 12087
rect 10318 12084 10324 12096
rect 10275 12056 10324 12084
rect 10275 12053 10287 12056
rect 10229 12047 10287 12053
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 13170 12084 13176 12096
rect 13131 12056 13176 12084
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13354 12084 13360 12096
rect 13315 12056 13360 12084
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 14200 12084 14228 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14826 12220 14832 12232
rect 14783 12192 14832 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 17402 12220 17408 12232
rect 17363 12192 17408 12220
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 14550 12112 14556 12164
rect 14608 12161 14614 12164
rect 14608 12155 14637 12161
rect 14625 12121 14637 12155
rect 14608 12115 14637 12121
rect 15648 12155 15706 12161
rect 15648 12121 15660 12155
rect 15694 12152 15706 12155
rect 17494 12152 17500 12164
rect 15694 12124 17500 12152
rect 15694 12121 15706 12124
rect 15648 12115 15706 12121
rect 14608 12112 14614 12115
rect 17494 12112 17500 12124
rect 17552 12112 17558 12164
rect 14826 12084 14832 12096
rect 14200 12056 14832 12084
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 17218 12084 17224 12096
rect 17179 12056 17224 12084
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 1104 11994 18860 12016
rect 1104 11942 6880 11994
rect 6932 11942 6944 11994
rect 6996 11942 7008 11994
rect 7060 11942 7072 11994
rect 7124 11942 7136 11994
rect 7188 11942 12811 11994
rect 12863 11942 12875 11994
rect 12927 11942 12939 11994
rect 12991 11942 13003 11994
rect 13055 11942 13067 11994
rect 13119 11942 18860 11994
rect 1104 11920 18860 11942
rect 6917 11883 6975 11889
rect 6917 11849 6929 11883
rect 6963 11880 6975 11883
rect 7282 11880 7288 11892
rect 6963 11852 7288 11880
rect 6963 11849 6975 11852
rect 6917 11843 6975 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 10502 11880 10508 11892
rect 10008 11852 10508 11880
rect 10008 11840 10014 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 13909 11883 13967 11889
rect 13909 11849 13921 11883
rect 13955 11880 13967 11883
rect 14550 11880 14556 11892
rect 13955 11852 14556 11880
rect 13955 11849 13967 11852
rect 13909 11843 13967 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 16117 11883 16175 11889
rect 16117 11849 16129 11883
rect 16163 11880 16175 11883
rect 16206 11880 16212 11892
rect 16163 11852 16212 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 5813 11815 5871 11821
rect 5813 11781 5825 11815
rect 5859 11812 5871 11815
rect 7098 11812 7104 11824
rect 5859 11784 7104 11812
rect 5859 11781 5871 11784
rect 5813 11775 5871 11781
rect 7098 11772 7104 11784
rect 7156 11772 7162 11824
rect 8662 11812 8668 11824
rect 7208 11784 8668 11812
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11744 4951 11747
rect 4982 11744 4988 11756
rect 4939 11716 4988 11744
rect 4939 11713 4951 11716
rect 4893 11707 4951 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 5534 11744 5540 11756
rect 5132 11716 5177 11744
rect 5495 11716 5540 11744
rect 5132 11704 5138 11716
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11744 5687 11747
rect 5902 11744 5908 11756
rect 5675 11716 5908 11744
rect 5675 11713 5687 11716
rect 5629 11707 5687 11713
rect 5902 11704 5908 11716
rect 5960 11744 5966 11756
rect 7208 11753 7236 11784
rect 8662 11772 8668 11784
rect 8720 11772 8726 11824
rect 9214 11772 9220 11824
rect 9272 11812 9278 11824
rect 9858 11812 9864 11824
rect 9272 11784 9720 11812
rect 9771 11784 9864 11812
rect 9272 11772 9278 11784
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 5960 11716 7205 11744
rect 5960 11704 5966 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 6270 11568 6276 11620
rect 6328 11608 6334 11620
rect 7300 11608 7328 11707
rect 7374 11704 7380 11756
rect 7432 11744 7438 11756
rect 7432 11716 7477 11744
rect 7432 11704 7438 11716
rect 7558 11704 7564 11756
rect 7616 11744 7622 11756
rect 8849 11747 8907 11753
rect 7616 11716 7661 11744
rect 7616 11704 7622 11716
rect 8849 11713 8861 11747
rect 8895 11744 8907 11747
rect 9030 11744 9036 11756
rect 8895 11716 9036 11744
rect 8895 11713 8907 11716
rect 8849 11707 8907 11713
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9582 11744 9588 11756
rect 9543 11716 9588 11744
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 9692 11753 9720 11784
rect 9858 11772 9864 11784
rect 9916 11812 9922 11824
rect 10226 11812 10232 11824
rect 9916 11784 10232 11812
rect 9916 11772 9922 11784
rect 10226 11772 10232 11784
rect 10284 11772 10290 11824
rect 15010 11821 15016 11824
rect 10781 11815 10839 11821
rect 10781 11812 10793 11815
rect 10428 11784 10793 11812
rect 9678 11747 9736 11753
rect 9678 11713 9690 11747
rect 9724 11713 9736 11747
rect 9950 11744 9956 11756
rect 9911 11716 9956 11744
rect 9678 11707 9736 11713
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 10091 11747 10149 11753
rect 10091 11713 10103 11747
rect 10137 11744 10149 11747
rect 10428 11744 10456 11784
rect 10781 11781 10793 11784
rect 10827 11781 10839 11815
rect 15004 11812 15016 11821
rect 14971 11784 15016 11812
rect 10781 11775 10839 11781
rect 15004 11775 15016 11784
rect 15010 11772 15016 11775
rect 15068 11772 15074 11824
rect 10137 11716 10456 11744
rect 10689 11747 10747 11753
rect 10137 11713 10149 11716
rect 10091 11707 10149 11713
rect 10689 11713 10701 11747
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 9125 11679 9183 11685
rect 9125 11645 9137 11679
rect 9171 11676 9183 11679
rect 10318 11676 10324 11688
rect 9171 11648 10324 11676
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 10318 11636 10324 11648
rect 10376 11676 10382 11688
rect 10704 11676 10732 11707
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 11664 11716 12081 11744
rect 11664 11704 11670 11716
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 12336 11747 12394 11753
rect 12336 11713 12348 11747
rect 12382 11744 12394 11747
rect 12710 11744 12716 11756
rect 12382 11716 12716 11744
rect 12382 11713 12394 11716
rect 12336 11707 12394 11713
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 14182 11744 14188 11756
rect 14139 11716 14188 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11744 14335 11747
rect 14550 11744 14556 11756
rect 14323 11716 14556 11744
rect 14323 11713 14335 11716
rect 14277 11707 14335 11713
rect 14550 11704 14556 11716
rect 14608 11704 14614 11756
rect 10376 11648 10732 11676
rect 10376 11636 10382 11648
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14734 11676 14740 11688
rect 14056 11648 14740 11676
rect 14056 11636 14062 11648
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 8018 11608 8024 11620
rect 6328 11580 8024 11608
rect 6328 11568 6334 11580
rect 8018 11568 8024 11580
rect 8076 11568 8082 11620
rect 9033 11611 9091 11617
rect 9033 11577 9045 11611
rect 9079 11608 9091 11611
rect 10134 11608 10140 11620
rect 9079 11580 10140 11608
rect 9079 11577 9091 11580
rect 9033 11571 9091 11577
rect 10134 11568 10140 11580
rect 10192 11568 10198 11620
rect 4430 11500 4436 11552
rect 4488 11540 4494 11552
rect 4893 11543 4951 11549
rect 4893 11540 4905 11543
rect 4488 11512 4905 11540
rect 4488 11500 4494 11512
rect 4893 11509 4905 11512
rect 4939 11509 4951 11543
rect 4893 11503 4951 11509
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5684 11512 5825 11540
rect 5684 11500 5690 11512
rect 5813 11509 5825 11512
rect 5859 11509 5871 11543
rect 5813 11503 5871 11509
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7926 11540 7932 11552
rect 7156 11512 7932 11540
rect 7156 11500 7162 11512
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8662 11540 8668 11552
rect 8623 11512 8668 11540
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 10229 11543 10287 11549
rect 10229 11509 10241 11543
rect 10275 11540 10287 11543
rect 11514 11540 11520 11552
rect 10275 11512 11520 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 13446 11540 13452 11552
rect 13407 11512 13452 11540
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 1104 11450 18860 11472
rect 1104 11398 3915 11450
rect 3967 11398 3979 11450
rect 4031 11398 4043 11450
rect 4095 11398 4107 11450
rect 4159 11398 4171 11450
rect 4223 11398 9846 11450
rect 9898 11398 9910 11450
rect 9962 11398 9974 11450
rect 10026 11398 10038 11450
rect 10090 11398 10102 11450
rect 10154 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 15904 11450
rect 15956 11398 15968 11450
rect 16020 11398 16032 11450
rect 16084 11398 18860 11450
rect 1104 11376 18860 11398
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7432 11308 7757 11336
rect 7432 11296 7438 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10376 11308 10517 11336
rect 10376 11296 10382 11308
rect 10505 11305 10517 11308
rect 10551 11305 10563 11339
rect 10505 11299 10563 11305
rect 11422 11296 11428 11348
rect 11480 11336 11486 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 11480 11308 11529 11336
rect 11480 11296 11486 11308
rect 11517 11305 11529 11308
rect 11563 11305 11575 11339
rect 11517 11299 11575 11305
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13722 11336 13728 11348
rect 13228 11308 13728 11336
rect 13228 11296 13234 11308
rect 13722 11296 13728 11308
rect 13780 11336 13786 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13780 11308 14105 11336
rect 13780 11296 13786 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14550 11336 14556 11348
rect 14511 11308 14556 11336
rect 14093 11299 14151 11305
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15654 11336 15660 11348
rect 15335 11308 15660 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 4982 11228 4988 11280
rect 5040 11268 5046 11280
rect 11701 11271 11759 11277
rect 5040 11240 7512 11268
rect 5040 11228 5046 11240
rect 6270 11200 6276 11212
rect 6231 11172 6276 11200
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 7374 11200 7380 11212
rect 6748 11172 7380 11200
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3844 11104 3985 11132
rect 3844 11092 3850 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11132 6239 11135
rect 6748 11132 6776 11172
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7484 11200 7512 11240
rect 11701 11237 11713 11271
rect 11747 11268 11759 11271
rect 15470 11268 15476 11280
rect 11747 11240 15476 11268
rect 11747 11237 11759 11240
rect 11701 11231 11759 11237
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 7650 11200 7656 11212
rect 7484 11172 7656 11200
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 8846 11160 8852 11212
rect 8904 11200 8910 11212
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 8904 11172 9137 11200
rect 8904 11160 8910 11172
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 12066 11200 12072 11212
rect 11204 11172 12072 11200
rect 11204 11160 11210 11172
rect 12066 11160 12072 11172
rect 12124 11200 12130 11212
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 12124 11172 12173 11200
rect 12124 11160 12130 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12161 11163 12219 11169
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 13538 11200 13544 11212
rect 12483 11172 13544 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 6227 11104 6776 11132
rect 6825 11135 6883 11141
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11132 7251 11135
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7239 11104 7849 11132
rect 7239 11101 7251 11104
rect 7193 11095 7251 11101
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 4246 11073 4252 11076
rect 4240 11064 4252 11073
rect 4207 11036 4252 11064
rect 4240 11027 4252 11036
rect 4246 11024 4252 11027
rect 4304 11024 4310 11076
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 6196 11064 6224 11095
rect 5132 11036 6224 11064
rect 5132 11024 5138 11036
rect 5368 11005 5396 11036
rect 5353 10999 5411 11005
rect 5353 10965 5365 10999
rect 5399 10965 5411 10999
rect 5810 10996 5816 11008
rect 5771 10968 5816 10996
rect 5353 10959 5411 10965
rect 5810 10956 5816 10968
rect 5868 10956 5874 11008
rect 6840 10996 6868 11095
rect 7024 11064 7052 11095
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 7984 11104 8029 11132
rect 7984 11092 7990 11104
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 9381 11135 9439 11141
rect 9381 11132 9393 11135
rect 8720 11104 9393 11132
rect 8720 11092 8726 11104
rect 9381 11101 9393 11104
rect 9427 11101 9439 11135
rect 9381 11095 9439 11101
rect 7282 11064 7288 11076
rect 7024 11036 7288 11064
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 11333 11067 11391 11073
rect 7432 11036 9352 11064
rect 7432 11024 7438 11036
rect 9324 11008 9352 11036
rect 11333 11033 11345 11067
rect 11379 11064 11391 11067
rect 12452 11064 12480 11163
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 14090 11160 14096 11212
rect 14148 11200 14154 11212
rect 14185 11203 14243 11209
rect 14185 11200 14197 11203
rect 14148 11172 14197 11200
rect 14148 11160 14154 11172
rect 14185 11169 14197 11172
rect 14231 11169 14243 11203
rect 14185 11163 14243 11169
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 13504 11104 14381 11132
rect 13504 11092 13510 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14734 11092 14740 11144
rect 14792 11132 14798 11144
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 14792 11104 16681 11132
rect 14792 11092 14798 11104
rect 16669 11101 16681 11104
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 11379 11036 12480 11064
rect 11379 11033 11391 11036
rect 11333 11027 11391 11033
rect 13354 11024 13360 11076
rect 13412 11064 13418 11076
rect 14093 11067 14151 11073
rect 14093 11064 14105 11067
rect 13412 11036 14105 11064
rect 13412 11024 13418 11036
rect 14093 11033 14105 11036
rect 14139 11033 14151 11067
rect 14093 11027 14151 11033
rect 16424 11067 16482 11073
rect 16424 11033 16436 11067
rect 16470 11064 16482 11067
rect 17218 11064 17224 11076
rect 16470 11036 17224 11064
rect 16470 11033 16482 11036
rect 16424 11027 16482 11033
rect 17218 11024 17224 11036
rect 17276 11024 17282 11076
rect 7742 10996 7748 11008
rect 6840 10968 7748 10996
rect 7742 10956 7748 10968
rect 7800 10956 7806 11008
rect 9306 10956 9312 11008
rect 9364 10956 9370 11008
rect 11514 10956 11520 11008
rect 11572 11005 11578 11008
rect 11572 10999 11591 11005
rect 11579 10965 11591 10999
rect 11572 10959 11591 10965
rect 11572 10956 11578 10959
rect 1104 10906 18860 10928
rect 1104 10854 6880 10906
rect 6932 10854 6944 10906
rect 6996 10854 7008 10906
rect 7060 10854 7072 10906
rect 7124 10854 7136 10906
rect 7188 10854 12811 10906
rect 12863 10854 12875 10906
rect 12927 10854 12939 10906
rect 12991 10854 13003 10906
rect 13055 10854 13067 10906
rect 13119 10854 18860 10906
rect 1104 10832 18860 10854
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 4246 10724 4252 10736
rect 4207 10696 4252 10724
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 4709 10727 4767 10733
rect 4709 10693 4721 10727
rect 4755 10724 4767 10727
rect 5184 10724 5212 10755
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 7984 10764 8401 10792
rect 7984 10752 7990 10764
rect 8389 10761 8401 10764
rect 8435 10761 8447 10795
rect 8389 10755 8447 10761
rect 8941 10795 8999 10801
rect 8941 10761 8953 10795
rect 8987 10792 8999 10795
rect 9582 10792 9588 10804
rect 8987 10764 9588 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 10468 10764 10609 10792
rect 10468 10752 10474 10764
rect 10597 10761 10609 10764
rect 10643 10792 10655 10795
rect 11422 10792 11428 10804
rect 10643 10764 11428 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 14001 10795 14059 10801
rect 14001 10761 14013 10795
rect 14047 10792 14059 10795
rect 14274 10792 14280 10804
rect 14047 10764 14280 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 14642 10792 14648 10804
rect 14603 10764 14648 10792
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 7650 10724 7656 10736
rect 4755 10696 5212 10724
rect 7611 10696 7656 10724
rect 4755 10693 4767 10696
rect 4709 10687 4767 10693
rect 7650 10684 7656 10696
rect 7708 10684 7714 10736
rect 7742 10684 7748 10736
rect 7800 10724 7806 10736
rect 7800 10696 8524 10724
rect 7800 10684 7806 10696
rect 4430 10656 4436 10668
rect 4391 10628 4436 10656
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 4798 10656 4804 10668
rect 4663 10628 4804 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 5810 10656 5816 10668
rect 5583 10628 5816 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 5960 10628 6561 10656
rect 5960 10616 5966 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 7668 10656 7696 10684
rect 8202 10656 8208 10668
rect 7668 10628 8208 10656
rect 6549 10619 6607 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8496 10665 8524 10696
rect 9306 10684 9312 10736
rect 9364 10724 9370 10736
rect 9766 10724 9772 10736
rect 9364 10696 9444 10724
rect 9364 10684 9370 10696
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10656 9183 10659
rect 9214 10656 9220 10668
rect 9171 10628 9220 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10557 4399 10591
rect 5626 10588 5632 10600
rect 5587 10560 5632 10588
rect 4341 10551 4399 10557
rect 4356 10520 4384 10551
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 6328 10560 6469 10588
rect 6328 10548 6334 10560
rect 6457 10557 6469 10560
rect 6503 10557 6515 10591
rect 8312 10588 8340 10619
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 9416 10665 9444 10696
rect 9508 10696 9772 10724
rect 9508 10665 9536 10696
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12161 10727 12219 10733
rect 12161 10724 12173 10727
rect 12124 10696 12173 10724
rect 12124 10684 12130 10696
rect 12161 10693 12173 10696
rect 12207 10693 12219 10727
rect 12161 10687 12219 10693
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9674 10656 9680 10668
rect 9635 10628 9680 10656
rect 9493 10619 9551 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 10318 10656 10324 10668
rect 10183 10628 10324 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 13170 10656 13176 10668
rect 13083 10628 13176 10656
rect 13170 10616 13176 10628
rect 13228 10656 13234 10668
rect 13538 10656 13544 10668
rect 13228 10628 13544 10656
rect 13228 10616 13234 10628
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 13814 10656 13820 10668
rect 13775 10628 13820 10656
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 14458 10656 14464 10668
rect 14419 10628 14464 10656
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 6457 10551 6515 10557
rect 7300 10560 8340 10588
rect 9309 10591 9367 10597
rect 7300 10532 7328 10560
rect 9309 10557 9321 10591
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 4614 10520 4620 10532
rect 4356 10492 4620 10520
rect 4614 10480 4620 10492
rect 4672 10520 4678 10532
rect 5994 10520 6000 10532
rect 4672 10492 6000 10520
rect 4672 10480 4678 10492
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 6917 10523 6975 10529
rect 6917 10489 6929 10523
rect 6963 10520 6975 10523
rect 7006 10520 7012 10532
rect 6963 10492 7012 10520
rect 6963 10489 6975 10492
rect 6917 10483 6975 10489
rect 7006 10480 7012 10492
rect 7064 10520 7070 10532
rect 7282 10520 7288 10532
rect 7064 10492 7288 10520
rect 7064 10480 7070 10492
rect 7282 10480 7288 10492
rect 7340 10480 7346 10532
rect 9324 10520 9352 10551
rect 10226 10548 10232 10600
rect 10284 10548 10290 10600
rect 10594 10548 10600 10600
rect 10652 10588 10658 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 10652 10560 12449 10588
rect 10652 10548 10658 10560
rect 12437 10557 12449 10560
rect 12483 10588 12495 10591
rect 12526 10588 12532 10600
rect 12483 10560 12532 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13722 10588 13728 10600
rect 13403 10560 13728 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 10244 10520 10272 10548
rect 9324 10492 10272 10520
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 7708 10424 7757 10452
rect 7708 10412 7714 10424
rect 7745 10421 7757 10424
rect 7791 10421 7803 10455
rect 7745 10415 7803 10421
rect 10413 10455 10471 10461
rect 10413 10421 10425 10455
rect 10459 10452 10471 10455
rect 10502 10452 10508 10464
rect 10459 10424 10508 10452
rect 10459 10421 10471 10424
rect 10413 10415 10471 10421
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 12894 10412 12900 10464
rect 12952 10452 12958 10464
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12952 10424 13001 10452
rect 12952 10412 12958 10424
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 12989 10415 13047 10421
rect 1104 10362 18860 10384
rect 1104 10310 3915 10362
rect 3967 10310 3979 10362
rect 4031 10310 4043 10362
rect 4095 10310 4107 10362
rect 4159 10310 4171 10362
rect 4223 10310 9846 10362
rect 9898 10310 9910 10362
rect 9962 10310 9974 10362
rect 10026 10310 10038 10362
rect 10090 10310 10102 10362
rect 10154 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 15904 10362
rect 15956 10310 15968 10362
rect 16020 10310 16032 10362
rect 16084 10310 18860 10362
rect 1104 10288 18860 10310
rect 5169 10251 5227 10257
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 5902 10248 5908 10260
rect 5215 10220 5908 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 7006 10248 7012 10260
rect 6104 10220 7012 10248
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 6104 10189 6132 10220
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 11790 10208 11796 10260
rect 11848 10248 11854 10260
rect 11885 10251 11943 10257
rect 11885 10248 11897 10251
rect 11848 10220 11897 10248
rect 11848 10208 11854 10220
rect 11885 10217 11897 10220
rect 11931 10217 11943 10251
rect 12710 10248 12716 10260
rect 12671 10220 12716 10248
rect 11885 10211 11943 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 5997 10183 6055 10189
rect 5997 10180 6009 10183
rect 5868 10152 6009 10180
rect 5868 10140 5874 10152
rect 5997 10149 6009 10152
rect 6043 10149 6055 10183
rect 5997 10143 6055 10149
rect 6089 10183 6147 10189
rect 6089 10149 6101 10183
rect 6135 10149 6147 10183
rect 6089 10143 6147 10149
rect 6917 10183 6975 10189
rect 6917 10149 6929 10183
rect 6963 10180 6975 10183
rect 7282 10180 7288 10192
rect 6963 10152 7288 10180
rect 6963 10149 6975 10152
rect 6917 10143 6975 10149
rect 7282 10140 7288 10152
rect 7340 10140 7346 10192
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5534 10112 5540 10124
rect 5399 10084 5540 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 6638 10112 6644 10124
rect 6328 10084 6644 10112
rect 6328 10072 6334 10084
rect 6638 10072 6644 10084
rect 6696 10112 6702 10124
rect 6825 10115 6883 10121
rect 6825 10112 6837 10115
rect 6696 10084 6837 10112
rect 6696 10072 6702 10084
rect 6825 10081 6837 10084
rect 6871 10112 6883 10115
rect 7650 10112 7656 10124
rect 6871 10084 7656 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7650 10072 7656 10084
rect 7708 10112 7714 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7708 10084 7849 10112
rect 7708 10072 7714 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 12158 10112 12164 10124
rect 11563 10084 12164 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 5074 10044 5080 10056
rect 5035 10016 5080 10044
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 7006 10044 7012 10056
rect 6967 10016 7012 10044
rect 6181 10007 6239 10013
rect 5353 9979 5411 9985
rect 5353 9945 5365 9979
rect 5399 9976 5411 9979
rect 5920 9976 5948 10007
rect 5399 9948 5948 9976
rect 6196 9976 6224 10007
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7929 10047 7987 10053
rect 7929 10044 7941 10047
rect 7147 10016 7941 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 7929 10013 7941 10016
rect 7975 10044 7987 10047
rect 8386 10044 8392 10056
rect 7975 10016 8392 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 11422 10044 11428 10056
rect 11383 10016 11428 10044
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 11606 10044 11612 10056
rect 11567 10016 11612 10044
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10044 11759 10047
rect 11974 10044 11980 10056
rect 11747 10016 11980 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 12894 10044 12900 10056
rect 12855 10016 12900 10044
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 7742 9976 7748 9988
rect 6196 9948 7748 9976
rect 5399 9945 5411 9948
rect 5353 9939 5411 9945
rect 7742 9936 7748 9948
rect 7800 9936 7806 9988
rect 6362 9908 6368 9920
rect 6323 9880 6368 9908
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 7432 9880 7573 9908
rect 7432 9868 7438 9880
rect 7561 9877 7573 9880
rect 7607 9877 7619 9911
rect 7561 9871 7619 9877
rect 1104 9818 18860 9840
rect 1104 9766 6880 9818
rect 6932 9766 6944 9818
rect 6996 9766 7008 9818
rect 7060 9766 7072 9818
rect 7124 9766 7136 9818
rect 7188 9766 12811 9818
rect 12863 9766 12875 9818
rect 12927 9766 12939 9818
rect 12991 9766 13003 9818
rect 13055 9766 13067 9818
rect 13119 9766 18860 9818
rect 1104 9744 18860 9766
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 17494 9704 17500 9716
rect 12584 9676 17500 9704
rect 12584 9664 12590 9676
rect 17494 9664 17500 9676
rect 17552 9704 17558 9716
rect 17862 9704 17868 9716
rect 17552 9676 17868 9704
rect 17552 9664 17558 9676
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 6457 9639 6515 9645
rect 6457 9636 6469 9639
rect 5592 9608 6469 9636
rect 5592 9596 5598 9608
rect 6457 9605 6469 9608
rect 6503 9605 6515 9639
rect 6638 9636 6644 9648
rect 6599 9608 6644 9636
rect 6457 9599 6515 9605
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 7742 9636 7748 9648
rect 6788 9608 7604 9636
rect 7703 9608 7748 9636
rect 6788 9596 6794 9608
rect 7576 9580 7604 9608
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 10502 9636 10508 9648
rect 7852 9608 10508 9636
rect 4982 9568 4988 9580
rect 4943 9540 4988 9568
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9537 5227 9571
rect 7282 9568 7288 9580
rect 7243 9540 7288 9568
rect 5169 9531 5227 9537
rect 5184 9500 5212 9531
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 7432 9540 7477 9568
rect 7432 9528 7438 9540
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 7616 9540 7709 9568
rect 7616 9528 7622 9540
rect 5258 9500 5264 9512
rect 5171 9472 5264 9500
rect 5258 9460 5264 9472
rect 5316 9500 5322 9512
rect 7852 9500 7880 9608
rect 10502 9596 10508 9608
rect 10560 9596 10566 9648
rect 8846 9528 8852 9580
rect 8904 9568 8910 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 8904 9540 9597 9568
rect 8904 9528 8910 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 9852 9571 9910 9577
rect 9852 9537 9864 9571
rect 9898 9568 9910 9571
rect 10226 9568 10232 9580
rect 9898 9540 10232 9568
rect 9898 9537 9910 9540
rect 9852 9531 9910 9537
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 5316 9472 7880 9500
rect 5316 9460 5322 9472
rect 7469 9435 7527 9441
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 7650 9432 7656 9444
rect 7515 9404 7656 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 7650 9392 7656 9404
rect 7708 9392 7714 9444
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 4985 9367 5043 9373
rect 4985 9364 4997 9367
rect 4764 9336 4997 9364
rect 4764 9324 4770 9336
rect 4985 9333 4997 9336
rect 5031 9333 5043 9367
rect 4985 9327 5043 9333
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10744 9336 10977 9364
rect 10744 9324 10750 9336
rect 10965 9333 10977 9336
rect 11011 9333 11023 9367
rect 10965 9327 11023 9333
rect 1104 9274 18860 9296
rect 1104 9222 3915 9274
rect 3967 9222 3979 9274
rect 4031 9222 4043 9274
rect 4095 9222 4107 9274
rect 4159 9222 4171 9274
rect 4223 9222 9846 9274
rect 9898 9222 9910 9274
rect 9962 9222 9974 9274
rect 10026 9222 10038 9274
rect 10090 9222 10102 9274
rect 10154 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 15904 9274
rect 15956 9222 15968 9274
rect 16020 9222 16032 9274
rect 16084 9222 18860 9274
rect 1104 9200 18860 9222
rect 4706 9160 4712 9172
rect 4667 9132 4712 9160
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 10226 9160 10232 9172
rect 10187 9132 10232 9160
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 11149 9163 11207 9169
rect 11149 9129 11161 9163
rect 11195 9160 11207 9163
rect 11422 9160 11428 9172
rect 11195 9132 11428 9160
rect 11195 9129 11207 9132
rect 11149 9123 11207 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 7561 9095 7619 9101
rect 7561 9061 7573 9095
rect 7607 9092 7619 9095
rect 8018 9092 8024 9104
rect 7607 9064 8024 9092
rect 7607 9061 7619 9064
rect 7561 9055 7619 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 4614 9024 4620 9036
rect 4575 8996 4620 9024
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 11425 9027 11483 9033
rect 11425 9024 11437 9027
rect 10560 8996 11437 9024
rect 10560 8984 10566 8996
rect 11425 8993 11437 8996
rect 11471 8993 11483 9027
rect 11425 8987 11483 8993
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 4798 8956 4804 8968
rect 4759 8928 4804 8956
rect 4798 8916 4804 8928
rect 4856 8956 4862 8968
rect 6546 8956 6552 8968
rect 4856 8928 6552 8956
rect 4856 8916 4862 8928
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 6779 8928 7389 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7377 8925 7389 8928
rect 7423 8956 7435 8959
rect 7834 8956 7840 8968
rect 7423 8928 7840 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 7834 8916 7840 8928
rect 7892 8956 7898 8968
rect 8202 8956 8208 8968
rect 7892 8928 8208 8956
rect 7892 8916 7898 8928
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 10410 8956 10416 8968
rect 10371 8928 10416 8956
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 10744 8928 11345 8956
rect 10744 8916 10750 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 11645 8959 11703 8965
rect 11572 8928 11617 8956
rect 11572 8916 11578 8928
rect 11645 8925 11657 8959
rect 11691 8956 11703 8959
rect 11882 8956 11888 8968
rect 11691 8928 11888 8956
rect 11691 8925 11703 8928
rect 11645 8919 11703 8925
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 4522 8888 4528 8900
rect 4483 8860 4528 8888
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 4982 8888 4988 8900
rect 4943 8860 4988 8888
rect 4982 8848 4988 8860
rect 5040 8848 5046 8900
rect 1104 8730 18860 8752
rect 1104 8678 6880 8730
rect 6932 8678 6944 8730
rect 6996 8678 7008 8730
rect 7060 8678 7072 8730
rect 7124 8678 7136 8730
rect 7188 8678 12811 8730
rect 12863 8678 12875 8730
rect 12927 8678 12939 8730
rect 12991 8678 13003 8730
rect 13055 8678 13067 8730
rect 13119 8678 18860 8730
rect 1104 8656 18860 8678
rect 5258 8616 5264 8628
rect 5219 8588 5264 8616
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 10410 8616 10416 8628
rect 10371 8588 10416 8616
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11974 8576 11980 8628
rect 12032 8616 12038 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 12032 8588 12081 8616
rect 12032 8576 12038 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 12069 8579 12127 8585
rect 4148 8551 4206 8557
rect 4148 8517 4160 8551
rect 4194 8548 4206 8551
rect 4522 8548 4528 8560
rect 4194 8520 4528 8548
rect 4194 8517 4206 8520
rect 4148 8511 4206 8517
rect 4522 8508 4528 8520
rect 4580 8508 4586 8560
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11164 8520 11713 8548
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 3881 8483 3939 8489
rect 3881 8480 3893 8483
rect 3844 8452 3893 8480
rect 3844 8440 3850 8452
rect 3881 8449 3893 8452
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 7432 8452 7757 8480
rect 7432 8440 7438 8452
rect 7745 8449 7757 8452
rect 7791 8480 7803 8483
rect 7834 8480 7840 8492
rect 7791 8452 7840 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 10962 8480 10968 8492
rect 10643 8452 10968 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 8018 8412 8024 8424
rect 7979 8384 8024 8412
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 10502 8372 10508 8424
rect 10560 8412 10566 8424
rect 10781 8415 10839 8421
rect 10781 8412 10793 8415
rect 10560 8384 10793 8412
rect 10560 8372 10566 8384
rect 10781 8381 10793 8384
rect 10827 8412 10839 8415
rect 11164 8412 11192 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 11701 8511 11759 8517
rect 11790 8480 11796 8492
rect 11751 8452 11796 8480
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 11974 8480 11980 8492
rect 11931 8452 11980 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 13170 8440 13176 8492
rect 13228 8480 13234 8492
rect 14277 8483 14335 8489
rect 14277 8480 14289 8483
rect 13228 8452 14289 8480
rect 13228 8440 13234 8452
rect 14277 8449 14289 8452
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 10827 8384 11192 8412
rect 14461 8415 14519 8421
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 14461 8381 14473 8415
rect 14507 8412 14519 8415
rect 14642 8412 14648 8424
rect 14507 8384 14648 8412
rect 14507 8381 14519 8384
rect 14461 8375 14519 8381
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 7926 8344 7932 8356
rect 7887 8316 7932 8344
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 10744 8316 11529 8344
rect 10744 8304 10750 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7800 8248 7849 8276
rect 7800 8236 7806 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 14090 8276 14096 8288
rect 14051 8248 14096 8276
rect 7837 8239 7895 8245
rect 14090 8236 14096 8248
rect 14148 8236 14154 8288
rect 1104 8186 18860 8208
rect 1104 8134 3915 8186
rect 3967 8134 3979 8186
rect 4031 8134 4043 8186
rect 4095 8134 4107 8186
rect 4159 8134 4171 8186
rect 4223 8134 9846 8186
rect 9898 8134 9910 8186
rect 9962 8134 9974 8186
rect 10026 8134 10038 8186
rect 10090 8134 10102 8186
rect 10154 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 15904 8186
rect 15956 8134 15968 8186
rect 16020 8134 16032 8186
rect 16084 8134 18860 8186
rect 1104 8112 18860 8134
rect 8018 8072 8024 8084
rect 7979 8044 8024 8072
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 14240 8044 14565 8072
rect 14240 8032 14246 8044
rect 14553 8041 14565 8044
rect 14599 8041 14611 8075
rect 14918 8072 14924 8084
rect 14879 8044 14924 8072
rect 14553 8035 14611 8041
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 8202 7936 8208 7948
rect 8163 7908 8208 7936
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 14921 7939 14979 7945
rect 14921 7905 14933 7939
rect 14967 7936 14979 7939
rect 15378 7936 15384 7948
rect 14967 7908 15384 7936
rect 14967 7905 14979 7908
rect 14921 7899 14979 7905
rect 15378 7896 15384 7908
rect 15436 7896 15442 7948
rect 7742 7868 7748 7880
rect 7703 7840 7748 7868
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 11793 7871 11851 7877
rect 7892 7840 7937 7868
rect 7892 7828 7898 7840
rect 11793 7837 11805 7871
rect 11839 7868 11851 7871
rect 12066 7868 12072 7880
rect 11839 7840 12072 7868
rect 11839 7837 11851 7840
rect 11793 7831 11851 7837
rect 12066 7828 12072 7840
rect 12124 7868 12130 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 12124 7840 12633 7868
rect 12124 7828 12130 7840
rect 12621 7837 12633 7840
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 14090 7868 14096 7880
rect 13403 7840 14096 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14734 7868 14740 7880
rect 14695 7840 14740 7868
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 14642 7760 14648 7812
rect 14700 7800 14706 7812
rect 15013 7803 15071 7809
rect 15013 7800 15025 7803
rect 14700 7772 15025 7800
rect 14700 7760 14706 7772
rect 15013 7769 15025 7772
rect 15059 7769 15071 7803
rect 15013 7763 15071 7769
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11609 7735 11667 7741
rect 11609 7732 11621 7735
rect 11112 7704 11621 7732
rect 11112 7692 11118 7704
rect 11609 7701 11621 7704
rect 11655 7701 11667 7735
rect 11609 7695 11667 7701
rect 12805 7735 12863 7741
rect 12805 7701 12817 7735
rect 12851 7732 12863 7735
rect 13354 7732 13360 7744
rect 12851 7704 13360 7732
rect 12851 7701 12863 7704
rect 12805 7695 12863 7701
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 13538 7732 13544 7744
rect 13499 7704 13544 7732
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 1104 7642 18860 7664
rect 1104 7590 6880 7642
rect 6932 7590 6944 7642
rect 6996 7590 7008 7642
rect 7060 7590 7072 7642
rect 7124 7590 7136 7642
rect 7188 7590 12811 7642
rect 12863 7590 12875 7642
rect 12927 7590 12939 7642
rect 12991 7590 13003 7642
rect 13055 7590 13067 7642
rect 13119 7590 18860 7642
rect 1104 7568 18860 7590
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 9493 7531 9551 7537
rect 9493 7528 9505 7531
rect 8536 7500 9505 7528
rect 8536 7488 8542 7500
rect 9493 7497 9505 7500
rect 9539 7497 9551 7531
rect 11514 7528 11520 7540
rect 11475 7500 11520 7528
rect 9493 7491 9551 7497
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 8846 7460 8852 7472
rect 8128 7432 8852 7460
rect 8128 7401 8156 7432
rect 8846 7420 8852 7432
rect 8904 7420 8910 7472
rect 13538 7420 13544 7472
rect 13596 7460 13602 7472
rect 14246 7463 14304 7469
rect 14246 7460 14258 7463
rect 13596 7432 14258 7460
rect 13596 7420 13602 7432
rect 14246 7429 14258 7432
rect 14292 7429 14304 7463
rect 14246 7423 14304 7429
rect 8386 7401 8392 7404
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8380 7355 8392 7401
rect 8444 7392 8450 7404
rect 10505 7395 10563 7401
rect 8444 7364 8480 7392
rect 8386 7352 8392 7355
rect 8444 7352 8450 7364
rect 10505 7361 10517 7395
rect 10551 7361 10563 7395
rect 10686 7392 10692 7404
rect 10647 7364 10692 7392
rect 10505 7355 10563 7361
rect 10520 7324 10548 7355
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 11882 7392 11888 7404
rect 11843 7364 11888 7392
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12618 7392 12624 7404
rect 12579 7364 12624 7392
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 11054 7324 11060 7336
rect 10520 7296 11060 7324
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11790 7324 11796 7336
rect 11751 7296 11796 7324
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 13998 7324 14004 7336
rect 13959 7296 14004 7324
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10321 7191 10379 7197
rect 10321 7188 10333 7191
rect 10284 7160 10333 7188
rect 10284 7148 10290 7160
rect 10321 7157 10333 7160
rect 10367 7157 10379 7191
rect 10321 7151 10379 7157
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 10928 7160 11897 7188
rect 10928 7148 10934 7160
rect 11885 7157 11897 7160
rect 11931 7188 11943 7191
rect 11974 7188 11980 7200
rect 11931 7160 11980 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 12434 7188 12440 7200
rect 12395 7160 12440 7188
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 15378 7188 15384 7200
rect 15291 7160 15384 7188
rect 15378 7148 15384 7160
rect 15436 7188 15442 7200
rect 16206 7188 16212 7200
rect 15436 7160 16212 7188
rect 15436 7148 15442 7160
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 1104 7098 18860 7120
rect 1104 7046 3915 7098
rect 3967 7046 3979 7098
rect 4031 7046 4043 7098
rect 4095 7046 4107 7098
rect 4159 7046 4171 7098
rect 4223 7046 9846 7098
rect 9898 7046 9910 7098
rect 9962 7046 9974 7098
rect 10026 7046 10038 7098
rect 10090 7046 10102 7098
rect 10154 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 15904 7098
rect 15956 7046 15968 7098
rect 16020 7046 16032 7098
rect 16084 7046 18860 7098
rect 1104 7024 18860 7046
rect 8297 6987 8355 6993
rect 8297 6953 8309 6987
rect 8343 6984 8355 6987
rect 8386 6984 8392 6996
rect 8343 6956 8392 6984
rect 8343 6953 8355 6956
rect 8297 6947 8355 6953
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 14921 6919 14979 6925
rect 14921 6916 14933 6919
rect 14792 6888 14933 6916
rect 14792 6876 14798 6888
rect 14921 6885 14933 6888
rect 14967 6885 14979 6919
rect 14921 6879 14979 6885
rect 15749 6919 15807 6925
rect 15749 6885 15761 6919
rect 15795 6914 15807 6919
rect 15795 6886 15829 6914
rect 15795 6885 15807 6886
rect 15749 6879 15807 6885
rect 8110 6848 8116 6860
rect 7944 6820 8116 6848
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 7524 6752 7665 6780
rect 7524 6740 7530 6752
rect 7653 6749 7665 6752
rect 7699 6749 7711 6783
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7653 6743 7711 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 7944 6789 7972 6820
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9490 6848 9496 6860
rect 8904 6820 9496 6848
rect 8904 6808 8910 6820
rect 9490 6808 9496 6820
rect 9548 6848 9554 6860
rect 11422 6848 11428 6860
rect 9548 6820 11428 6848
rect 9548 6808 9554 6820
rect 11422 6808 11428 6820
rect 11480 6848 11486 6860
rect 11885 6851 11943 6857
rect 11885 6848 11897 6851
rect 11480 6820 11897 6848
rect 11480 6808 11486 6820
rect 11885 6817 11897 6820
rect 11931 6817 11943 6851
rect 11885 6811 11943 6817
rect 14369 6851 14427 6857
rect 14369 6817 14381 6851
rect 14415 6848 14427 6851
rect 14826 6848 14832 6860
rect 14415 6820 14832 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 15764 6848 15792 6879
rect 15068 6820 15792 6848
rect 15068 6808 15074 6820
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8478 6780 8484 6792
rect 8067 6752 8484 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 10226 6780 10232 6792
rect 10187 6752 10232 6780
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 12152 6783 12210 6789
rect 12152 6749 12164 6783
rect 12198 6780 12210 6783
rect 12434 6780 12440 6792
rect 12198 6752 12440 6780
rect 12198 6749 12210 6752
rect 12152 6743 12210 6749
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 15102 6780 15108 6792
rect 14056 6752 15108 6780
rect 14056 6740 14062 6752
rect 15102 6740 15108 6752
rect 15160 6780 15166 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 15160 6752 17141 6780
rect 15160 6740 15166 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 14366 6672 14372 6724
rect 14424 6712 14430 6724
rect 14737 6715 14795 6721
rect 14737 6712 14749 6715
rect 14424 6684 14749 6712
rect 14424 6672 14430 6684
rect 14737 6681 14749 6684
rect 14783 6712 14795 6715
rect 14918 6712 14924 6724
rect 14783 6684 14924 6712
rect 14783 6681 14795 6684
rect 14737 6675 14795 6681
rect 14918 6672 14924 6684
rect 14976 6672 14982 6724
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 16862 6715 16920 6721
rect 16862 6712 16874 6715
rect 16816 6684 16874 6712
rect 16816 6672 16822 6684
rect 16862 6681 16874 6684
rect 16908 6681 16920 6715
rect 16862 6675 16920 6681
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10045 6647 10103 6653
rect 10045 6644 10057 6647
rect 9824 6616 10057 6644
rect 9824 6604 9830 6616
rect 10045 6613 10057 6616
rect 10091 6613 10103 6647
rect 10045 6607 10103 6613
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 12492 6616 13277 6644
rect 12492 6604 12498 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 14550 6644 14556 6656
rect 14511 6616 14556 6644
rect 13265 6607 13323 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 14645 6647 14703 6653
rect 14645 6613 14657 6647
rect 14691 6644 14703 6647
rect 16206 6644 16212 6656
rect 14691 6616 16212 6644
rect 14691 6613 14703 6616
rect 14645 6607 14703 6613
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 1104 6554 18860 6576
rect 1104 6502 6880 6554
rect 6932 6502 6944 6554
rect 6996 6502 7008 6554
rect 7060 6502 7072 6554
rect 7124 6502 7136 6554
rect 7188 6502 12811 6554
rect 12863 6502 12875 6554
rect 12927 6502 12939 6554
rect 12991 6502 13003 6554
rect 13055 6502 13067 6554
rect 13119 6502 18860 6554
rect 1104 6480 18860 6502
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7800 6412 7849 6440
rect 7800 6400 7806 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 11664 6412 12173 6440
rect 11664 6400 11670 6412
rect 12161 6409 12173 6412
rect 12207 6409 12219 6443
rect 12434 6440 12440 6452
rect 12395 6412 12440 6440
rect 12161 6403 12219 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 12676 6412 13185 6440
rect 12676 6400 12682 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 14001 6443 14059 6449
rect 14001 6409 14013 6443
rect 14047 6440 14059 6443
rect 14550 6440 14556 6452
rect 14047 6412 14556 6440
rect 14047 6409 14059 6412
rect 14001 6403 14059 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 15102 6400 15108 6452
rect 15160 6400 15166 6452
rect 6546 6332 6552 6384
rect 6604 6372 6610 6384
rect 15120 6372 15148 6400
rect 6604 6344 7144 6372
rect 6604 6332 6610 6344
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6304 4951 6307
rect 5258 6304 5264 6316
rect 4939 6276 5264 6304
rect 4939 6273 4951 6276
rect 4893 6267 4951 6273
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 7116 6313 7144 6344
rect 12360 6344 13492 6372
rect 15120 6344 15424 6372
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 6788 6276 6929 6304
rect 6788 6264 6794 6276
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6273 7159 6307
rect 7558 6304 7564 6316
rect 7519 6276 7564 6304
rect 7101 6267 7159 6273
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 7650 6264 7656 6316
rect 7708 6304 7714 6316
rect 7708 6276 7753 6304
rect 7708 6264 7714 6276
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12360 6313 12388 6344
rect 12345 6307 12403 6313
rect 12345 6304 12357 6307
rect 12216 6276 12357 6304
rect 12216 6264 12222 6276
rect 12345 6273 12357 6276
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6304 12587 6307
rect 12618 6304 12624 6316
rect 12575 6276 12624 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 13354 6304 13360 6316
rect 13315 6276 13360 6304
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 13464 6313 13492 6344
rect 15396 6313 15424 6344
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 15125 6307 15183 6313
rect 15125 6273 15137 6307
rect 15171 6304 15183 6307
rect 15381 6307 15439 6313
rect 15171 6276 15332 6304
rect 15171 6273 15183 6276
rect 15125 6267 15183 6273
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6236 5043 6239
rect 5534 6236 5540 6248
rect 5031 6208 5540 6236
rect 5031 6205 5043 6208
rect 4985 6199 5043 6205
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8110 6236 8116 6248
rect 7883 6208 8116 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 15304 6236 15332 6276
rect 15381 6273 15393 6307
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 15562 6264 15568 6316
rect 15620 6304 15626 6316
rect 16025 6307 16083 6313
rect 16025 6304 16037 6307
rect 15620 6276 16037 6304
rect 15620 6264 15626 6276
rect 16025 6273 16037 6276
rect 16071 6273 16083 6307
rect 17310 6304 17316 6316
rect 17271 6276 17316 6304
rect 16025 6267 16083 6273
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17494 6304 17500 6316
rect 17455 6276 17500 6304
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 15304 6208 15884 6236
rect 12250 6128 12256 6180
rect 12308 6168 12314 6180
rect 15856 6177 15884 6208
rect 12713 6171 12771 6177
rect 12713 6168 12725 6171
rect 12308 6140 12725 6168
rect 12308 6128 12314 6140
rect 12713 6137 12725 6140
rect 12759 6137 12771 6171
rect 12713 6131 12771 6137
rect 15841 6171 15899 6177
rect 15841 6137 15853 6171
rect 15887 6137 15899 6171
rect 15841 6131 15899 6137
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 7009 6103 7067 6109
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7466 6100 7472 6112
rect 7055 6072 7472 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 17129 6103 17187 6109
rect 17129 6100 17141 6103
rect 17000 6072 17141 6100
rect 17000 6060 17006 6072
rect 17129 6069 17141 6072
rect 17175 6069 17187 6103
rect 17129 6063 17187 6069
rect 1104 6010 18860 6032
rect 1104 5958 3915 6010
rect 3967 5958 3979 6010
rect 4031 5958 4043 6010
rect 4095 5958 4107 6010
rect 4159 5958 4171 6010
rect 4223 5958 9846 6010
rect 9898 5958 9910 6010
rect 9962 5958 9974 6010
rect 10026 5958 10038 6010
rect 10090 5958 10102 6010
rect 10154 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 15904 6010
rect 15956 5958 15968 6010
rect 16020 5958 16032 6010
rect 16084 5958 18860 6010
rect 1104 5936 18860 5958
rect 4801 5899 4859 5905
rect 4801 5865 4813 5899
rect 4847 5896 4859 5899
rect 4982 5896 4988 5908
rect 4847 5868 4988 5896
rect 4847 5865 4859 5868
rect 4801 5859 4859 5865
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 6730 5896 6736 5908
rect 6691 5868 6736 5896
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 10870 5896 10876 5908
rect 10831 5868 10876 5896
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 12161 5899 12219 5905
rect 12161 5896 12173 5899
rect 11940 5868 12173 5896
rect 11940 5856 11946 5868
rect 12161 5865 12173 5868
rect 12207 5865 12219 5899
rect 12618 5896 12624 5908
rect 12579 5868 12624 5896
rect 12161 5859 12219 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 15473 5899 15531 5905
rect 15473 5865 15485 5899
rect 15519 5896 15531 5899
rect 15562 5896 15568 5908
rect 15519 5868 15568 5896
rect 15519 5865 15531 5868
rect 15473 5859 15531 5865
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 16758 5896 16764 5908
rect 16719 5868 16764 5896
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 17957 5899 18015 5905
rect 17957 5896 17969 5899
rect 17368 5868 17969 5896
rect 17368 5856 17374 5868
rect 17957 5865 17969 5868
rect 18003 5865 18015 5899
rect 17957 5859 18015 5865
rect 6638 5788 6644 5840
rect 6696 5828 6702 5840
rect 9214 5828 9220 5840
rect 6696 5800 9220 5828
rect 6696 5788 6702 5800
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 12636 5828 12664 5856
rect 11348 5800 12664 5828
rect 4522 5720 4528 5772
rect 4580 5760 4586 5772
rect 4985 5763 5043 5769
rect 4985 5760 4997 5763
rect 4580 5732 4997 5760
rect 4580 5720 4586 5732
rect 4985 5729 4997 5732
rect 5031 5729 5043 5763
rect 4985 5723 5043 5729
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 7650 5760 7656 5772
rect 7147 5732 7656 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 9490 5760 9496 5772
rect 9451 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 11348 5769 11376 5800
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5729 11391 5763
rect 12434 5760 12440 5772
rect 12395 5732 12440 5760
rect 11333 5723 11391 5729
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 14734 5720 14740 5772
rect 14792 5760 14798 5772
rect 15105 5763 15163 5769
rect 15105 5760 15117 5763
rect 14792 5732 15117 5760
rect 14792 5720 14798 5732
rect 15105 5729 15117 5732
rect 15151 5729 15163 5763
rect 15105 5723 15163 5729
rect 5074 5692 5080 5704
rect 5035 5664 5080 5692
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5592 5664 5917 5692
rect 5592 5652 5598 5664
rect 5905 5661 5917 5664
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5692 6147 5695
rect 6638 5692 6644 5704
rect 6135 5664 6644 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 5920 5624 5948 5655
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5692 7067 5695
rect 7558 5692 7564 5704
rect 7055 5664 7564 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8294 5692 8300 5704
rect 8255 5664 8300 5692
rect 8113 5655 8171 5661
rect 6730 5624 6736 5636
rect 5920 5596 6736 5624
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 7282 5584 7288 5636
rect 7340 5624 7346 5636
rect 7742 5624 7748 5636
rect 7340 5596 7748 5624
rect 7340 5584 7346 5596
rect 7742 5584 7748 5596
rect 7800 5624 7806 5636
rect 8128 5624 8156 5655
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 9766 5701 9772 5704
rect 9760 5692 9772 5701
rect 9727 5664 9772 5692
rect 9760 5655 9772 5664
rect 9766 5652 9772 5655
rect 9824 5652 9830 5704
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11112 5664 11529 5692
rect 11112 5652 11118 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 12345 5695 12403 5701
rect 12345 5692 12357 5695
rect 12308 5664 12357 5692
rect 12308 5652 12314 5664
rect 12345 5661 12357 5664
rect 12391 5692 12403 5695
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 12391 5664 13093 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5692 13323 5695
rect 13354 5692 13360 5704
rect 13311 5664 13360 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 13354 5652 13360 5664
rect 13412 5652 13418 5704
rect 14366 5692 14372 5704
rect 14327 5664 14372 5692
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14507 5664 15301 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 15289 5661 15301 5664
rect 15335 5692 15347 5695
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15335 5664 16129 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 7800 5596 8156 5624
rect 11701 5627 11759 5633
rect 7800 5584 7806 5596
rect 11701 5593 11713 5627
rect 11747 5593 11759 5627
rect 11701 5587 11759 5593
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 5997 5559 6055 5565
rect 5997 5556 6009 5559
rect 5592 5528 6009 5556
rect 5592 5516 5598 5528
rect 5997 5525 6009 5528
rect 6043 5525 6055 5559
rect 8110 5556 8116 5568
rect 8071 5528 8116 5556
rect 5997 5519 6055 5525
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 11716 5556 11744 5587
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 12621 5627 12679 5633
rect 12621 5624 12633 5627
rect 12216 5596 12633 5624
rect 12216 5584 12222 5596
rect 12621 5593 12633 5596
rect 12667 5593 12679 5627
rect 13372 5624 13400 5652
rect 14476 5624 14504 5655
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 16942 5692 16948 5704
rect 16264 5664 16309 5692
rect 16903 5664 16948 5692
rect 16264 5652 16270 5664
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 17862 5652 17868 5704
rect 17920 5692 17926 5704
rect 18141 5695 18199 5701
rect 18141 5692 18153 5695
rect 17920 5664 18153 5692
rect 17920 5652 17926 5664
rect 18141 5661 18153 5664
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 13372 5596 14504 5624
rect 12621 5587 12679 5593
rect 13354 5556 13360 5568
rect 11716 5528 13360 5556
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 14274 5556 14280 5568
rect 13495 5528 14280 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 14645 5559 14703 5565
rect 14645 5525 14657 5559
rect 14691 5556 14703 5559
rect 14918 5556 14924 5568
rect 14691 5528 14924 5556
rect 14691 5525 14703 5528
rect 14645 5519 14703 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 15933 5559 15991 5565
rect 15933 5556 15945 5559
rect 15620 5528 15945 5556
rect 15620 5516 15626 5528
rect 15933 5525 15945 5528
rect 15979 5525 15991 5559
rect 15933 5519 15991 5525
rect 1104 5466 18860 5488
rect 1104 5414 6880 5466
rect 6932 5414 6944 5466
rect 6996 5414 7008 5466
rect 7060 5414 7072 5466
rect 7124 5414 7136 5466
rect 7188 5414 12811 5466
rect 12863 5414 12875 5466
rect 12927 5414 12939 5466
rect 12991 5414 13003 5466
rect 13055 5414 13067 5466
rect 13119 5414 18860 5466
rect 1104 5392 18860 5414
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 5132 5324 5273 5352
rect 5132 5312 5138 5324
rect 5261 5321 5273 5324
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 8294 5312 8300 5364
rect 8352 5312 8358 5364
rect 12158 5352 12164 5364
rect 12119 5324 12164 5352
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 15381 5355 15439 5361
rect 15381 5352 15393 5355
rect 14792 5324 15393 5352
rect 14792 5312 14798 5324
rect 15381 5321 15393 5324
rect 15427 5321 15439 5355
rect 15381 5315 15439 5321
rect 6365 5287 6423 5293
rect 6365 5284 6377 5287
rect 4632 5256 6377 5284
rect 4632 5225 4660 5256
rect 6365 5253 6377 5256
rect 6411 5253 6423 5287
rect 6730 5284 6736 5296
rect 6691 5256 6736 5284
rect 6365 5247 6423 5253
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 7374 5284 7380 5296
rect 7300 5256 7380 5284
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 5537 5219 5595 5225
rect 4847 5188 5304 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 5276 5157 5304 5188
rect 5537 5185 5549 5219
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6638 5216 6644 5228
rect 6595 5188 6644 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5442 5148 5448 5160
rect 5307 5120 5448 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 4709 5083 4767 5089
rect 4709 5049 4721 5083
rect 4755 5080 4767 5083
rect 5350 5080 5356 5092
rect 4755 5052 5356 5080
rect 4755 5049 4767 5052
rect 4709 5043 4767 5049
rect 5350 5040 5356 5052
rect 5408 5080 5414 5092
rect 5552 5080 5580 5179
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 7300 5225 7328 5256
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 8018 5284 8024 5296
rect 7576 5256 8024 5284
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 7285 5179 7343 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7576 5225 7604 5256
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 8312 5284 8340 5312
rect 8757 5287 8815 5293
rect 8757 5284 8769 5287
rect 8312 5256 8769 5284
rect 8757 5253 8769 5256
rect 8803 5253 8815 5287
rect 8757 5247 8815 5253
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 7742 5216 7748 5228
rect 7699 5188 7748 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 8352 5188 8585 5216
rect 8352 5176 8358 5188
rect 8573 5185 8585 5188
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 9999 5188 10425 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 10870 5216 10876 5228
rect 10827 5188 10876 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 10612 5148 10640 5179
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11514 5216 11520 5228
rect 11475 5188 11520 5216
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 13285 5219 13343 5225
rect 13285 5185 13297 5219
rect 13331 5216 13343 5219
rect 13446 5216 13452 5228
rect 13331 5188 13452 5216
rect 13331 5185 13343 5188
rect 13285 5179 13343 5185
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5216 13599 5219
rect 13998 5216 14004 5228
rect 13587 5188 14004 5216
rect 13587 5185 13599 5188
rect 13541 5179 13599 5185
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 14268 5219 14326 5225
rect 14268 5185 14280 5219
rect 14314 5216 14326 5219
rect 14734 5216 14740 5228
rect 14314 5188 14740 5216
rect 14314 5185 14326 5188
rect 14268 5179 14326 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 11054 5148 11060 5160
rect 10612 5120 11060 5148
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 5408 5052 5580 5080
rect 5408 5040 5414 5052
rect 5445 5015 5503 5021
rect 5445 4981 5457 5015
rect 5491 5012 5503 5015
rect 5534 5012 5540 5024
rect 5491 4984 5540 5012
rect 5491 4981 5503 4984
rect 5445 4975 5503 4981
rect 5534 4972 5540 4984
rect 5592 5012 5598 5024
rect 6362 5012 6368 5024
rect 5592 4984 6368 5012
rect 5592 4972 5598 4984
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 7558 4972 7564 5024
rect 7616 5012 7622 5024
rect 7929 5015 7987 5021
rect 7929 5012 7941 5015
rect 7616 4984 7941 5012
rect 7616 4972 7622 4984
rect 7929 4981 7941 4984
rect 7975 4981 7987 5015
rect 8386 5012 8392 5024
rect 8347 4984 8392 5012
rect 7929 4975 7987 4981
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9732 4984 9781 5012
rect 9732 4972 9738 4984
rect 9769 4981 9781 4984
rect 9815 4981 9827 5015
rect 11698 5012 11704 5024
rect 11659 4984 11704 5012
rect 9769 4975 9827 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 1104 4922 18860 4944
rect 1104 4870 3915 4922
rect 3967 4870 3979 4922
rect 4031 4870 4043 4922
rect 4095 4870 4107 4922
rect 4159 4870 4171 4922
rect 4223 4870 9846 4922
rect 9898 4870 9910 4922
rect 9962 4870 9974 4922
rect 10026 4870 10038 4922
rect 10090 4870 10102 4922
rect 10154 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 15904 4922
rect 15956 4870 15968 4922
rect 16020 4870 16032 4922
rect 16084 4870 18860 4922
rect 1104 4848 18860 4870
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7650 4808 7656 4820
rect 7607 4780 7656 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 7800 4780 8217 4808
rect 7800 4768 7806 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 10965 4811 11023 4817
rect 10965 4777 10977 4811
rect 11011 4808 11023 4811
rect 11146 4808 11152 4820
rect 11011 4780 11152 4808
rect 11011 4777 11023 4780
rect 10965 4771 11023 4777
rect 11146 4768 11152 4780
rect 11204 4808 11210 4820
rect 11790 4808 11796 4820
rect 11204 4780 11796 4808
rect 11204 4768 11210 4780
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12676 4780 12817 4808
rect 12676 4768 12682 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 12805 4771 12863 4777
rect 13446 4768 13452 4820
rect 13504 4808 13510 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13504 4780 14105 4808
rect 13504 4768 13510 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14734 4808 14740 4820
rect 14695 4780 14740 4808
rect 14093 4771 14151 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 6638 4740 6644 4752
rect 6472 4712 6644 4740
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4672 5503 4675
rect 5534 4672 5540 4684
rect 5491 4644 5540 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6472 4613 6500 4712
rect 6638 4700 6644 4712
rect 6696 4740 6702 4752
rect 7466 4740 7472 4752
rect 6696 4712 7472 4740
rect 6696 4700 6702 4712
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 8110 4672 8116 4684
rect 7484 4644 8116 4672
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6546 4604 6604 4610
rect 6546 4570 6558 4604
rect 6592 4570 6604 4604
rect 6546 4564 6604 4570
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 6825 4607 6883 4613
rect 6696 4576 6741 4604
rect 6696 4564 6702 4576
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 7374 4604 7380 4616
rect 6871 4576 7380 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 7484 4613 7512 4644
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 9585 4675 9643 4681
rect 9585 4672 9597 4675
rect 9548 4644 9597 4672
rect 9548 4632 9554 4644
rect 9585 4641 9597 4644
rect 9631 4641 9643 4675
rect 11422 4672 11428 4684
rect 11383 4644 11428 4672
rect 9585 4635 9643 4641
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 8386 4604 8392 4616
rect 7699 4576 8392 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 11698 4613 11704 4616
rect 9841 4607 9899 4613
rect 9841 4604 9853 4607
rect 9732 4576 9853 4604
rect 9732 4564 9738 4576
rect 9841 4573 9853 4576
rect 9887 4573 9899 4607
rect 11692 4604 11704 4613
rect 11659 4576 11704 4604
rect 9841 4567 9899 4573
rect 11692 4567 11704 4576
rect 11698 4564 11704 4567
rect 11756 4564 11762 4616
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 13412 4576 13461 4604
rect 13412 4564 13418 4576
rect 13449 4573 13461 4576
rect 13495 4573 13507 4607
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 13449 4567 13507 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14918 4604 14924 4616
rect 14879 4576 14924 4604
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 15562 4604 15568 4616
rect 15523 4576 15568 4604
rect 15562 4564 15568 4576
rect 15620 4564 15626 4616
rect 6564 4536 6592 4564
rect 8294 4536 8300 4548
rect 6564 4508 6684 4536
rect 8255 4508 8300 4536
rect 5718 4468 5724 4480
rect 5679 4440 5724 4468
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 6178 4468 6184 4480
rect 6139 4440 6184 4468
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 6656 4468 6684 4508
rect 8294 4496 8300 4508
rect 8352 4496 8358 4548
rect 13262 4468 13268 4480
rect 6604 4440 6684 4468
rect 13223 4440 13268 4468
rect 6604 4428 6610 4440
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 15378 4468 15384 4480
rect 15339 4440 15384 4468
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 1104 4378 18860 4400
rect 1104 4326 6880 4378
rect 6932 4326 6944 4378
rect 6996 4326 7008 4378
rect 7060 4326 7072 4378
rect 7124 4326 7136 4378
rect 7188 4326 12811 4378
rect 12863 4326 12875 4378
rect 12927 4326 12939 4378
rect 12991 4326 13003 4378
rect 13055 4326 13067 4378
rect 13119 4326 18860 4378
rect 1104 4304 18860 4326
rect 6549 4267 6607 4273
rect 6549 4233 6561 4267
rect 6595 4264 6607 4267
rect 6638 4264 6644 4276
rect 6595 4236 6644 4264
rect 6595 4233 6607 4236
rect 6549 4227 6607 4233
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8665 4267 8723 4273
rect 8665 4264 8677 4267
rect 8352 4236 8677 4264
rect 8352 4224 8358 4236
rect 8665 4233 8677 4236
rect 8711 4233 8723 4267
rect 10502 4264 10508 4276
rect 10463 4236 10508 4264
rect 8665 4227 8723 4233
rect 10502 4224 10508 4236
rect 10560 4224 10566 4276
rect 9490 4196 9496 4208
rect 7392 4168 7696 4196
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5776 4100 6377 4128
rect 5776 4088 5782 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6546 4128 6552 4140
rect 6507 4100 6552 4128
rect 6365 4091 6423 4097
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 7392 4128 7420 4168
rect 7558 4137 7564 4140
rect 7552 4128 7564 4137
rect 7331 4100 7420 4128
rect 7519 4100 7564 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 7552 4091 7564 4100
rect 6086 4020 6092 4072
rect 6144 4060 6150 4072
rect 7300 4060 7328 4091
rect 7558 4088 7564 4091
rect 7616 4088 7622 4140
rect 7668 4128 7696 4168
rect 9140 4168 9496 4196
rect 9140 4137 9168 4168
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 12836 4199 12894 4205
rect 12836 4165 12848 4199
rect 12882 4196 12894 4199
rect 13262 4196 13268 4208
rect 12882 4168 13268 4196
rect 12882 4165 12894 4168
rect 12836 4159 12894 4165
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 15378 4196 15384 4208
rect 14936 4168 15384 4196
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 7668 4100 9137 4128
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9392 4131 9450 4137
rect 9392 4097 9404 4131
rect 9438 4128 9450 4131
rect 9766 4128 9772 4140
rect 9438 4100 9772 4128
rect 9438 4097 9450 4100
rect 9392 4091 9450 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13998 4128 14004 4140
rect 13127 4100 14004 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 14849 4131 14907 4137
rect 14849 4097 14861 4131
rect 14895 4128 14907 4131
rect 14936 4128 14964 4168
rect 15378 4156 15384 4168
rect 15436 4156 15442 4208
rect 15102 4128 15108 4140
rect 14895 4100 14964 4128
rect 15063 4100 15108 4128
rect 14895 4097 14907 4100
rect 14849 4091 14907 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 15565 4131 15623 4137
rect 15565 4128 15577 4131
rect 15528 4100 15577 4128
rect 15528 4088 15534 4100
rect 15565 4097 15577 4100
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 6144 4032 7328 4060
rect 6144 4020 6150 4032
rect 13722 3992 13728 4004
rect 13683 3964 13728 3992
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 12158 3924 12164 3936
rect 11747 3896 12164 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 15749 3927 15807 3933
rect 15749 3893 15761 3927
rect 15795 3924 15807 3927
rect 16850 3924 16856 3936
rect 15795 3896 16856 3924
rect 15795 3893 15807 3896
rect 15749 3887 15807 3893
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 1104 3834 18860 3856
rect 1104 3782 3915 3834
rect 3967 3782 3979 3834
rect 4031 3782 4043 3834
rect 4095 3782 4107 3834
rect 4159 3782 4171 3834
rect 4223 3782 9846 3834
rect 9898 3782 9910 3834
rect 9962 3782 9974 3834
rect 10026 3782 10038 3834
rect 10090 3782 10102 3834
rect 10154 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 15904 3834
rect 15956 3782 15968 3834
rect 16020 3782 16032 3834
rect 16084 3782 18860 3834
rect 1104 3760 18860 3782
rect 7466 3720 7472 3732
rect 7427 3692 7472 3720
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 9766 3720 9772 3732
rect 9727 3692 9772 3720
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 11241 3723 11299 3729
rect 11241 3689 11253 3723
rect 11287 3720 11299 3723
rect 11514 3720 11520 3732
rect 11287 3692 11520 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 12526 3652 12532 3664
rect 8956 3624 12532 3652
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 8956 3593 8984 3624
rect 12526 3612 12532 3624
rect 12584 3612 12590 3664
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 11146 3584 11152 3596
rect 10919 3556 11152 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 6178 3476 6184 3528
rect 6236 3516 6242 3528
rect 6345 3519 6403 3525
rect 6345 3516 6357 3519
rect 6236 3488 6357 3516
rect 6236 3476 6242 3488
rect 6345 3485 6357 3488
rect 6391 3485 6403 3519
rect 9122 3516 9128 3528
rect 9083 3488 9128 3516
rect 6345 3479 6403 3485
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9355 3488 9965 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 11054 3516 11060 3528
rect 11015 3488 11060 3516
rect 9953 3479 10011 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 1104 3290 18860 3312
rect 1104 3238 6880 3290
rect 6932 3238 6944 3290
rect 6996 3238 7008 3290
rect 7060 3238 7072 3290
rect 7124 3238 7136 3290
rect 7188 3238 12811 3290
rect 12863 3238 12875 3290
rect 12927 3238 12939 3290
rect 12991 3238 13003 3290
rect 13055 3238 13067 3290
rect 13119 3238 18860 3290
rect 1104 3216 18860 3238
rect 1104 2746 18860 2768
rect 1104 2694 3915 2746
rect 3967 2694 3979 2746
rect 4031 2694 4043 2746
rect 4095 2694 4107 2746
rect 4159 2694 4171 2746
rect 4223 2694 9846 2746
rect 9898 2694 9910 2746
rect 9962 2694 9974 2746
rect 10026 2694 10038 2746
rect 10090 2694 10102 2746
rect 10154 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 15904 2746
rect 15956 2694 15968 2746
rect 16020 2694 16032 2746
rect 16084 2694 18860 2746
rect 1104 2672 18860 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 9122 2632 9128 2644
rect 1627 2604 9128 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8444 2400 8953 2428
rect 8444 2388 8450 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 16850 2428 16856 2440
rect 16811 2400 16856 2428
rect 8941 2391 8999 2397
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 1104 2202 18860 2224
rect 1104 2150 6880 2202
rect 6932 2150 6944 2202
rect 6996 2150 7008 2202
rect 7060 2150 7072 2202
rect 7124 2150 7136 2202
rect 7188 2150 12811 2202
rect 12863 2150 12875 2202
rect 12927 2150 12939 2202
rect 12991 2150 13003 2202
rect 13055 2150 13067 2202
rect 13119 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 3915 47302 3967 47354
rect 3979 47302 4031 47354
rect 4043 47302 4095 47354
rect 4107 47302 4159 47354
rect 4171 47302 4223 47354
rect 9846 47302 9898 47354
rect 9910 47302 9962 47354
rect 9974 47302 10026 47354
rect 10038 47302 10090 47354
rect 10102 47302 10154 47354
rect 15776 47302 15828 47354
rect 15840 47302 15892 47354
rect 15904 47302 15956 47354
rect 15968 47302 16020 47354
rect 16032 47302 16084 47354
rect 11060 47200 11112 47252
rect 19340 47200 19392 47252
rect 2780 47039 2832 47048
rect 2780 47005 2789 47039
rect 2789 47005 2823 47039
rect 2823 47005 2832 47039
rect 2780 46996 2832 47005
rect 17868 47039 17920 47048
rect 17868 47005 17877 47039
rect 17877 47005 17911 47039
rect 17911 47005 17920 47039
rect 17868 46996 17920 47005
rect 3240 46928 3292 46980
rect 6880 46758 6932 46810
rect 6944 46758 6996 46810
rect 7008 46758 7060 46810
rect 7072 46758 7124 46810
rect 7136 46758 7188 46810
rect 12811 46758 12863 46810
rect 12875 46758 12927 46810
rect 12939 46758 12991 46810
rect 13003 46758 13055 46810
rect 13067 46758 13119 46810
rect 3915 46214 3967 46266
rect 3979 46214 4031 46266
rect 4043 46214 4095 46266
rect 4107 46214 4159 46266
rect 4171 46214 4223 46266
rect 9846 46214 9898 46266
rect 9910 46214 9962 46266
rect 9974 46214 10026 46266
rect 10038 46214 10090 46266
rect 10102 46214 10154 46266
rect 15776 46214 15828 46266
rect 15840 46214 15892 46266
rect 15904 46214 15956 46266
rect 15968 46214 16020 46266
rect 16032 46214 16084 46266
rect 8852 45908 8904 45960
rect 9128 45951 9180 45960
rect 9128 45917 9137 45951
rect 9137 45917 9171 45951
rect 9171 45917 9180 45951
rect 9128 45908 9180 45917
rect 9220 45772 9272 45824
rect 6880 45670 6932 45722
rect 6944 45670 6996 45722
rect 7008 45670 7060 45722
rect 7072 45670 7124 45722
rect 7136 45670 7188 45722
rect 12811 45670 12863 45722
rect 12875 45670 12927 45722
rect 12939 45670 12991 45722
rect 13003 45670 13055 45722
rect 13067 45670 13119 45722
rect 6184 45364 6236 45416
rect 7932 45364 7984 45416
rect 8116 45364 8168 45416
rect 8852 45500 8904 45552
rect 8852 45296 8904 45348
rect 10324 45500 10376 45552
rect 10416 45432 10468 45484
rect 11520 45475 11572 45484
rect 11520 45441 11529 45475
rect 11529 45441 11563 45475
rect 11563 45441 11572 45475
rect 11520 45432 11572 45441
rect 12072 45432 12124 45484
rect 6920 45271 6972 45280
rect 6920 45237 6929 45271
rect 6929 45237 6963 45271
rect 6963 45237 6972 45271
rect 7472 45271 7524 45280
rect 6920 45228 6972 45237
rect 7472 45237 7481 45271
rect 7481 45237 7515 45271
rect 7515 45237 7524 45271
rect 7472 45228 7524 45237
rect 8668 45228 8720 45280
rect 9036 45228 9088 45280
rect 10232 45228 10284 45280
rect 13268 45228 13320 45280
rect 3915 45126 3967 45178
rect 3979 45126 4031 45178
rect 4043 45126 4095 45178
rect 4107 45126 4159 45178
rect 4171 45126 4223 45178
rect 9846 45126 9898 45178
rect 9910 45126 9962 45178
rect 9974 45126 10026 45178
rect 10038 45126 10090 45178
rect 10102 45126 10154 45178
rect 15776 45126 15828 45178
rect 15840 45126 15892 45178
rect 15904 45126 15956 45178
rect 15968 45126 16020 45178
rect 16032 45126 16084 45178
rect 6920 45024 6972 45076
rect 7380 45067 7432 45076
rect 7380 45033 7389 45067
rect 7389 45033 7423 45067
rect 7423 45033 7432 45067
rect 7380 45024 7432 45033
rect 17868 44956 17920 45008
rect 6368 44820 6420 44872
rect 7564 44863 7616 44872
rect 7564 44829 7573 44863
rect 7573 44829 7607 44863
rect 7607 44829 7616 44863
rect 7564 44820 7616 44829
rect 5816 44795 5868 44804
rect 5816 44761 5850 44795
rect 5850 44761 5868 44795
rect 8024 44820 8076 44872
rect 8300 44820 8352 44872
rect 8944 44863 8996 44872
rect 8944 44829 8953 44863
rect 8953 44829 8987 44863
rect 8987 44829 8996 44863
rect 8944 44820 8996 44829
rect 9036 44820 9088 44872
rect 10876 44863 10928 44872
rect 10876 44829 10885 44863
rect 10885 44829 10919 44863
rect 10919 44829 10928 44863
rect 10876 44820 10928 44829
rect 11428 44863 11480 44872
rect 5816 44752 5868 44761
rect 6552 44684 6604 44736
rect 10416 44752 10468 44804
rect 11428 44829 11437 44863
rect 11437 44829 11471 44863
rect 11471 44829 11480 44863
rect 11428 44820 11480 44829
rect 11612 44863 11664 44872
rect 11612 44829 11621 44863
rect 11621 44829 11655 44863
rect 11655 44829 11664 44863
rect 11612 44820 11664 44829
rect 12072 44863 12124 44872
rect 12072 44829 12081 44863
rect 12081 44829 12115 44863
rect 12115 44829 12124 44863
rect 12072 44820 12124 44829
rect 11336 44752 11388 44804
rect 8392 44684 8444 44736
rect 10324 44727 10376 44736
rect 10324 44693 10333 44727
rect 10333 44693 10367 44727
rect 10367 44693 10376 44727
rect 10324 44684 10376 44693
rect 10876 44684 10928 44736
rect 6880 44582 6932 44634
rect 6944 44582 6996 44634
rect 7008 44582 7060 44634
rect 7072 44582 7124 44634
rect 7136 44582 7188 44634
rect 12811 44582 12863 44634
rect 12875 44582 12927 44634
rect 12939 44582 12991 44634
rect 13003 44582 13055 44634
rect 13067 44582 13119 44634
rect 5816 44480 5868 44532
rect 7932 44480 7984 44532
rect 12072 44480 12124 44532
rect 1860 44387 1912 44396
rect 1860 44353 1869 44387
rect 1869 44353 1903 44387
rect 1903 44353 1912 44387
rect 1860 44344 1912 44353
rect 7380 44412 7432 44464
rect 7472 44455 7524 44464
rect 7472 44421 7490 44455
rect 7490 44421 7524 44455
rect 7472 44412 7524 44421
rect 5816 44387 5868 44396
rect 5816 44353 5825 44387
rect 5825 44353 5859 44387
rect 5859 44353 5868 44387
rect 5816 44344 5868 44353
rect 7840 44344 7892 44396
rect 8392 44387 8444 44396
rect 8392 44353 8401 44387
rect 8401 44353 8435 44387
rect 8435 44353 8444 44387
rect 8392 44344 8444 44353
rect 8668 44387 8720 44396
rect 8668 44353 8677 44387
rect 8677 44353 8711 44387
rect 8711 44353 8720 44387
rect 8668 44344 8720 44353
rect 10324 44344 10376 44396
rect 12808 44344 12860 44396
rect 13820 44344 13872 44396
rect 7748 44319 7800 44328
rect 7748 44285 7757 44319
rect 7757 44285 7791 44319
rect 7791 44285 7800 44319
rect 7748 44276 7800 44285
rect 8116 44208 8168 44260
rect 7472 44140 7524 44192
rect 9772 44140 9824 44192
rect 3915 44038 3967 44090
rect 3979 44038 4031 44090
rect 4043 44038 4095 44090
rect 4107 44038 4159 44090
rect 4171 44038 4223 44090
rect 9846 44038 9898 44090
rect 9910 44038 9962 44090
rect 9974 44038 10026 44090
rect 10038 44038 10090 44090
rect 10102 44038 10154 44090
rect 15776 44038 15828 44090
rect 15840 44038 15892 44090
rect 15904 44038 15956 44090
rect 15968 44038 16020 44090
rect 16032 44038 16084 44090
rect 5816 43936 5868 43988
rect 6460 43868 6512 43920
rect 7564 43936 7616 43988
rect 8668 43936 8720 43988
rect 10232 43936 10284 43988
rect 11428 43936 11480 43988
rect 12808 43936 12860 43988
rect 11612 43868 11664 43920
rect 13268 43911 13320 43920
rect 6184 43843 6236 43852
rect 6184 43809 6193 43843
rect 6193 43809 6227 43843
rect 6227 43809 6236 43843
rect 6184 43800 6236 43809
rect 6368 43732 6420 43784
rect 6552 43732 6604 43784
rect 10876 43800 10928 43852
rect 12256 43843 12308 43852
rect 12256 43809 12265 43843
rect 12265 43809 12299 43843
rect 12299 43809 12308 43843
rect 12256 43800 12308 43809
rect 13268 43877 13277 43911
rect 13277 43877 13311 43911
rect 13311 43877 13320 43911
rect 13268 43868 13320 43877
rect 7472 43732 7524 43784
rect 7748 43732 7800 43784
rect 8944 43775 8996 43784
rect 8944 43741 8953 43775
rect 8953 43741 8987 43775
rect 8987 43741 8996 43775
rect 8944 43732 8996 43741
rect 9220 43775 9272 43784
rect 9220 43741 9254 43775
rect 9254 43741 9272 43775
rect 10784 43775 10836 43784
rect 9220 43732 9272 43741
rect 10784 43741 10793 43775
rect 10793 43741 10827 43775
rect 10827 43741 10836 43775
rect 10784 43732 10836 43741
rect 11336 43775 11388 43784
rect 10232 43664 10284 43716
rect 10968 43596 11020 43648
rect 11336 43741 11345 43775
rect 11345 43741 11379 43775
rect 11379 43741 11388 43775
rect 11336 43732 11388 43741
rect 12440 43664 12492 43716
rect 11980 43639 12032 43648
rect 11980 43605 11989 43639
rect 11989 43605 12023 43639
rect 12023 43605 12032 43639
rect 11980 43596 12032 43605
rect 12532 43596 12584 43648
rect 13268 43596 13320 43648
rect 6880 43494 6932 43546
rect 6944 43494 6996 43546
rect 7008 43494 7060 43546
rect 7072 43494 7124 43546
rect 7136 43494 7188 43546
rect 12811 43494 12863 43546
rect 12875 43494 12927 43546
rect 12939 43494 12991 43546
rect 13003 43494 13055 43546
rect 13067 43494 13119 43546
rect 6460 43392 6512 43444
rect 10784 43392 10836 43444
rect 12440 43435 12492 43444
rect 12440 43401 12449 43435
rect 12449 43401 12483 43435
rect 12483 43401 12492 43435
rect 12440 43392 12492 43401
rect 7932 43324 7984 43376
rect 8576 43324 8628 43376
rect 10324 43367 10376 43376
rect 8116 43299 8168 43308
rect 8116 43265 8125 43299
rect 8125 43265 8159 43299
rect 8159 43265 8168 43299
rect 8116 43256 8168 43265
rect 8668 43256 8720 43308
rect 9220 43299 9272 43308
rect 9220 43265 9229 43299
rect 9229 43265 9263 43299
rect 9263 43265 9272 43299
rect 9220 43256 9272 43265
rect 9680 43299 9732 43308
rect 9680 43265 9694 43299
rect 9694 43265 9728 43299
rect 9728 43265 9732 43299
rect 10324 43333 10333 43367
rect 10333 43333 10367 43367
rect 10367 43333 10376 43367
rect 10324 43324 10376 43333
rect 10968 43324 11020 43376
rect 9680 43256 9732 43265
rect 10232 43188 10284 43240
rect 10784 43299 10836 43308
rect 10784 43265 10793 43299
rect 10793 43265 10827 43299
rect 10827 43265 10836 43299
rect 10784 43256 10836 43265
rect 11888 43256 11940 43308
rect 11980 43231 12032 43240
rect 9588 43120 9640 43172
rect 6552 43052 6604 43104
rect 7748 43052 7800 43104
rect 8300 43052 8352 43104
rect 10508 43095 10560 43104
rect 10508 43061 10517 43095
rect 10517 43061 10551 43095
rect 10551 43061 10560 43095
rect 10508 43052 10560 43061
rect 11980 43197 11989 43231
rect 11989 43197 12023 43231
rect 12023 43197 12032 43231
rect 11980 43188 12032 43197
rect 12532 43120 12584 43172
rect 10876 43052 10928 43104
rect 11612 43052 11664 43104
rect 3915 42950 3967 43002
rect 3979 42950 4031 43002
rect 4043 42950 4095 43002
rect 4107 42950 4159 43002
rect 4171 42950 4223 43002
rect 9846 42950 9898 43002
rect 9910 42950 9962 43002
rect 9974 42950 10026 43002
rect 10038 42950 10090 43002
rect 10102 42950 10154 43002
rect 15776 42950 15828 43002
rect 15840 42950 15892 43002
rect 15904 42950 15956 43002
rect 15968 42950 16020 43002
rect 16032 42950 16084 43002
rect 8300 42848 8352 42900
rect 6184 42780 6236 42832
rect 9036 42712 9088 42764
rect 10968 42755 11020 42764
rect 10968 42721 10977 42755
rect 10977 42721 11011 42755
rect 11011 42721 11020 42755
rect 10968 42712 11020 42721
rect 9680 42644 9732 42696
rect 9772 42644 9824 42696
rect 12440 42644 12492 42696
rect 9128 42508 9180 42560
rect 9588 42508 9640 42560
rect 6880 42406 6932 42458
rect 6944 42406 6996 42458
rect 7008 42406 7060 42458
rect 7072 42406 7124 42458
rect 7136 42406 7188 42458
rect 12811 42406 12863 42458
rect 12875 42406 12927 42458
rect 12939 42406 12991 42458
rect 13003 42406 13055 42458
rect 13067 42406 13119 42458
rect 9220 42304 9272 42356
rect 10508 42304 10560 42356
rect 8668 42236 8720 42288
rect 7656 42168 7708 42220
rect 7840 42168 7892 42220
rect 8392 42211 8444 42220
rect 8392 42177 8401 42211
rect 8401 42177 8435 42211
rect 8435 42177 8444 42211
rect 8392 42168 8444 42177
rect 8576 42211 8628 42220
rect 8576 42177 8585 42211
rect 8585 42177 8619 42211
rect 8619 42177 8628 42211
rect 8576 42168 8628 42177
rect 9588 42168 9640 42220
rect 9772 42168 9824 42220
rect 10876 42168 10928 42220
rect 11520 42168 11572 42220
rect 8484 42100 8536 42152
rect 7932 41964 7984 42016
rect 3915 41862 3967 41914
rect 3979 41862 4031 41914
rect 4043 41862 4095 41914
rect 4107 41862 4159 41914
rect 4171 41862 4223 41914
rect 9846 41862 9898 41914
rect 9910 41862 9962 41914
rect 9974 41862 10026 41914
rect 10038 41862 10090 41914
rect 10102 41862 10154 41914
rect 15776 41862 15828 41914
rect 15840 41862 15892 41914
rect 15904 41862 15956 41914
rect 15968 41862 16020 41914
rect 16032 41862 16084 41914
rect 6880 41318 6932 41370
rect 6944 41318 6996 41370
rect 7008 41318 7060 41370
rect 7072 41318 7124 41370
rect 7136 41318 7188 41370
rect 12811 41318 12863 41370
rect 12875 41318 12927 41370
rect 12939 41318 12991 41370
rect 13003 41318 13055 41370
rect 13067 41318 13119 41370
rect 8392 41216 8444 41268
rect 8300 41191 8352 41200
rect 8300 41157 8309 41191
rect 8309 41157 8343 41191
rect 8343 41157 8352 41191
rect 8300 41148 8352 41157
rect 8116 41123 8168 41132
rect 8116 41089 8125 41123
rect 8125 41089 8159 41123
rect 8159 41089 8168 41123
rect 8116 41080 8168 41089
rect 8392 41123 8444 41132
rect 8392 41089 8401 41123
rect 8401 41089 8435 41123
rect 8435 41089 8444 41123
rect 8392 41080 8444 41089
rect 8576 41080 8628 41132
rect 14464 41055 14516 41064
rect 14464 41021 14473 41055
rect 14473 41021 14507 41055
rect 14507 41021 14516 41055
rect 14464 41012 14516 41021
rect 16672 41080 16724 41132
rect 18144 41123 18196 41132
rect 18144 41089 18153 41123
rect 18153 41089 18187 41123
rect 18187 41089 18196 41123
rect 18144 41080 18196 41089
rect 15384 41012 15436 41064
rect 15476 40919 15528 40928
rect 15476 40885 15485 40919
rect 15485 40885 15519 40919
rect 15519 40885 15528 40919
rect 15476 40876 15528 40885
rect 16120 40919 16172 40928
rect 16120 40885 16129 40919
rect 16129 40885 16163 40919
rect 16163 40885 16172 40919
rect 16120 40876 16172 40885
rect 17960 40919 18012 40928
rect 17960 40885 17969 40919
rect 17969 40885 18003 40919
rect 18003 40885 18012 40919
rect 17960 40876 18012 40885
rect 3915 40774 3967 40826
rect 3979 40774 4031 40826
rect 4043 40774 4095 40826
rect 4107 40774 4159 40826
rect 4171 40774 4223 40826
rect 9846 40774 9898 40826
rect 9910 40774 9962 40826
rect 9974 40774 10026 40826
rect 10038 40774 10090 40826
rect 10102 40774 10154 40826
rect 15776 40774 15828 40826
rect 15840 40774 15892 40826
rect 15904 40774 15956 40826
rect 15968 40774 16020 40826
rect 16032 40774 16084 40826
rect 6644 40672 6696 40724
rect 8300 40715 8352 40724
rect 8300 40681 8309 40715
rect 8309 40681 8343 40715
rect 8343 40681 8352 40715
rect 8300 40672 8352 40681
rect 8392 40672 8444 40724
rect 6736 40400 6788 40452
rect 7748 40468 7800 40520
rect 9680 40468 9732 40520
rect 12624 40468 12676 40520
rect 14740 40468 14792 40520
rect 16120 40468 16172 40520
rect 6460 40332 6512 40384
rect 8300 40400 8352 40452
rect 15476 40400 15528 40452
rect 7932 40332 7984 40384
rect 12716 40332 12768 40384
rect 14648 40332 14700 40384
rect 17408 40375 17460 40384
rect 17408 40341 17417 40375
rect 17417 40341 17451 40375
rect 17451 40341 17460 40375
rect 17408 40332 17460 40341
rect 6880 40230 6932 40282
rect 6944 40230 6996 40282
rect 7008 40230 7060 40282
rect 7072 40230 7124 40282
rect 7136 40230 7188 40282
rect 12811 40230 12863 40282
rect 12875 40230 12927 40282
rect 12939 40230 12991 40282
rect 13003 40230 13055 40282
rect 13067 40230 13119 40282
rect 8116 40128 8168 40180
rect 8024 40060 8076 40112
rect 5632 40035 5684 40044
rect 5632 40001 5641 40035
rect 5641 40001 5675 40035
rect 5675 40001 5684 40035
rect 5632 39992 5684 40001
rect 6552 40035 6604 40044
rect 6552 40001 6561 40035
rect 6561 40001 6595 40035
rect 6595 40001 6604 40035
rect 6552 39992 6604 40001
rect 6644 39992 6696 40044
rect 7748 40035 7800 40044
rect 7748 40001 7766 40035
rect 7766 40001 7800 40035
rect 7748 39992 7800 40001
rect 7932 40035 7984 40044
rect 7932 40001 7941 40035
rect 7941 40001 7975 40035
rect 7975 40001 7984 40035
rect 7932 39992 7984 40001
rect 8760 40060 8812 40112
rect 12716 40060 12768 40112
rect 15384 40060 15436 40112
rect 8944 39992 8996 40044
rect 10232 39992 10284 40044
rect 12072 39992 12124 40044
rect 12532 39992 12584 40044
rect 15568 39992 15620 40044
rect 6000 39924 6052 39976
rect 6736 39924 6788 39976
rect 6828 39967 6880 39976
rect 6828 39933 6837 39967
rect 6837 39933 6871 39967
rect 6871 39933 6880 39967
rect 6828 39924 6880 39933
rect 10324 39924 10376 39976
rect 5540 39788 5592 39840
rect 5908 39788 5960 39840
rect 8116 39788 8168 39840
rect 10784 39831 10836 39840
rect 10784 39797 10793 39831
rect 10793 39797 10827 39831
rect 10827 39797 10836 39831
rect 10784 39788 10836 39797
rect 11704 39788 11756 39840
rect 13820 39924 13872 39976
rect 14740 39967 14792 39976
rect 14740 39933 14749 39967
rect 14749 39933 14783 39967
rect 14783 39933 14792 39967
rect 14740 39924 14792 39933
rect 16672 39967 16724 39976
rect 16672 39933 16681 39967
rect 16681 39933 16715 39967
rect 16715 39933 16724 39967
rect 16672 39924 16724 39933
rect 16120 39899 16172 39908
rect 16120 39865 16129 39899
rect 16129 39865 16163 39899
rect 16163 39865 16172 39899
rect 16120 39856 16172 39865
rect 13820 39788 13872 39840
rect 14464 39788 14516 39840
rect 15108 39788 15160 39840
rect 3915 39686 3967 39738
rect 3979 39686 4031 39738
rect 4043 39686 4095 39738
rect 4107 39686 4159 39738
rect 4171 39686 4223 39738
rect 9846 39686 9898 39738
rect 9910 39686 9962 39738
rect 9974 39686 10026 39738
rect 10038 39686 10090 39738
rect 10102 39686 10154 39738
rect 15776 39686 15828 39738
rect 15840 39686 15892 39738
rect 15904 39686 15956 39738
rect 15968 39686 16020 39738
rect 16032 39686 16084 39738
rect 9680 39584 9732 39636
rect 11888 39627 11940 39636
rect 11888 39593 11897 39627
rect 11897 39593 11931 39627
rect 11931 39593 11940 39627
rect 11888 39584 11940 39593
rect 12624 39584 12676 39636
rect 15108 39584 15160 39636
rect 15384 39584 15436 39636
rect 7564 39516 7616 39568
rect 10232 39559 10284 39568
rect 10232 39525 10241 39559
rect 10241 39525 10275 39559
rect 10275 39525 10284 39559
rect 10232 39516 10284 39525
rect 7380 39448 7432 39500
rect 9956 39491 10008 39500
rect 9956 39457 9965 39491
rect 9965 39457 9999 39491
rect 9999 39457 10008 39491
rect 9956 39448 10008 39457
rect 11060 39516 11112 39568
rect 12256 39516 12308 39568
rect 12532 39448 12584 39500
rect 3608 39380 3660 39432
rect 6368 39380 6420 39432
rect 8116 39423 8168 39432
rect 5908 39312 5960 39364
rect 6828 39312 6880 39364
rect 5724 39244 5776 39296
rect 8116 39389 8125 39423
rect 8125 39389 8159 39423
rect 8159 39389 8168 39423
rect 8116 39380 8168 39389
rect 11704 39423 11756 39432
rect 7932 39312 7984 39364
rect 9772 39312 9824 39364
rect 11704 39389 11713 39423
rect 11713 39389 11747 39423
rect 11747 39389 11756 39423
rect 11704 39380 11756 39389
rect 11796 39423 11848 39432
rect 11796 39389 11805 39423
rect 11805 39389 11839 39423
rect 11839 39389 11848 39423
rect 15200 39448 15252 39500
rect 11796 39380 11848 39389
rect 13452 39312 13504 39364
rect 14188 39312 14240 39364
rect 14648 39380 14700 39432
rect 15752 39516 15804 39568
rect 15660 39423 15712 39432
rect 15660 39389 15669 39423
rect 15669 39389 15703 39423
rect 15703 39389 15712 39423
rect 15660 39380 15712 39389
rect 17960 39312 18012 39364
rect 8484 39244 8536 39296
rect 10416 39244 10468 39296
rect 13176 39244 13228 39296
rect 14924 39287 14976 39296
rect 14924 39253 14933 39287
rect 14933 39253 14967 39287
rect 14967 39253 14976 39287
rect 14924 39244 14976 39253
rect 15936 39244 15988 39296
rect 6880 39142 6932 39194
rect 6944 39142 6996 39194
rect 7008 39142 7060 39194
rect 7072 39142 7124 39194
rect 7136 39142 7188 39194
rect 12811 39142 12863 39194
rect 12875 39142 12927 39194
rect 12939 39142 12991 39194
rect 13003 39142 13055 39194
rect 13067 39142 13119 39194
rect 6552 39040 6604 39092
rect 7932 39040 7984 39092
rect 8944 39083 8996 39092
rect 8944 39049 8953 39083
rect 8953 39049 8987 39083
rect 8987 39049 8996 39083
rect 8944 39040 8996 39049
rect 6368 38972 6420 39024
rect 7288 38972 7340 39024
rect 11060 39040 11112 39092
rect 12072 39083 12124 39092
rect 12072 39049 12081 39083
rect 12081 39049 12115 39083
rect 12115 39049 12124 39083
rect 12072 39040 12124 39049
rect 15108 39083 15160 39092
rect 15108 39049 15117 39083
rect 15117 39049 15151 39083
rect 15151 39049 15160 39083
rect 15108 39040 15160 39049
rect 15568 39040 15620 39092
rect 3608 38947 3660 38956
rect 3608 38913 3617 38947
rect 3617 38913 3651 38947
rect 3651 38913 3660 38947
rect 3608 38904 3660 38913
rect 3700 38904 3752 38956
rect 5724 38947 5776 38956
rect 5724 38913 5733 38947
rect 5733 38913 5767 38947
rect 5767 38913 5776 38947
rect 5724 38904 5776 38913
rect 6000 38904 6052 38956
rect 6644 38947 6696 38956
rect 6644 38913 6678 38947
rect 6678 38913 6696 38947
rect 8208 38947 8260 38956
rect 6644 38904 6696 38913
rect 8208 38913 8217 38947
rect 8217 38913 8251 38947
rect 8251 38913 8260 38947
rect 8208 38904 8260 38913
rect 8392 38947 8444 38956
rect 8392 38913 8401 38947
rect 8401 38913 8435 38947
rect 8435 38913 8444 38947
rect 8392 38904 8444 38913
rect 8760 38947 8812 38956
rect 8760 38913 8769 38947
rect 8769 38913 8803 38947
rect 8803 38913 8812 38947
rect 8760 38904 8812 38913
rect 10508 38972 10560 39024
rect 12440 38972 12492 39024
rect 9680 38947 9732 38956
rect 9680 38913 9689 38947
rect 9689 38913 9723 38947
rect 9723 38913 9732 38947
rect 10416 38947 10468 38956
rect 9680 38904 9732 38913
rect 10416 38913 10425 38947
rect 10425 38913 10459 38947
rect 10459 38913 10468 38947
rect 10416 38904 10468 38913
rect 6368 38879 6420 38888
rect 4528 38700 4580 38752
rect 6368 38845 6377 38879
rect 6377 38845 6411 38879
rect 6411 38845 6420 38879
rect 6368 38836 6420 38845
rect 8024 38836 8076 38888
rect 10232 38836 10284 38888
rect 10324 38768 10376 38820
rect 10600 38811 10652 38820
rect 10600 38777 10609 38811
rect 10609 38777 10643 38811
rect 10643 38777 10652 38811
rect 10600 38768 10652 38777
rect 12256 38904 12308 38956
rect 13820 38972 13872 39024
rect 14648 38972 14700 39024
rect 15660 38972 15712 39024
rect 13176 38947 13228 38956
rect 13176 38913 13210 38947
rect 13210 38913 13228 38947
rect 13176 38904 13228 38913
rect 14188 38904 14240 38956
rect 15200 38904 15252 38956
rect 15752 38904 15804 38956
rect 15936 38947 15988 38956
rect 15936 38913 15945 38947
rect 15945 38913 15979 38947
rect 15979 38913 15988 38947
rect 15936 38904 15988 38913
rect 11796 38836 11848 38888
rect 10968 38768 11020 38820
rect 7840 38700 7892 38752
rect 14188 38700 14240 38752
rect 14372 38700 14424 38752
rect 3915 38598 3967 38650
rect 3979 38598 4031 38650
rect 4043 38598 4095 38650
rect 4107 38598 4159 38650
rect 4171 38598 4223 38650
rect 9846 38598 9898 38650
rect 9910 38598 9962 38650
rect 9974 38598 10026 38650
rect 10038 38598 10090 38650
rect 10102 38598 10154 38650
rect 15776 38598 15828 38650
rect 15840 38598 15892 38650
rect 15904 38598 15956 38650
rect 15968 38598 16020 38650
rect 16032 38598 16084 38650
rect 12532 38539 12584 38548
rect 12532 38505 12541 38539
rect 12541 38505 12575 38539
rect 12575 38505 12584 38539
rect 12532 38496 12584 38505
rect 15200 38496 15252 38548
rect 6736 38428 6788 38480
rect 11060 38428 11112 38480
rect 8116 38360 8168 38412
rect 9772 38403 9824 38412
rect 9772 38369 9781 38403
rect 9781 38369 9815 38403
rect 9815 38369 9824 38403
rect 9772 38360 9824 38369
rect 10324 38360 10376 38412
rect 3792 38335 3844 38344
rect 3792 38301 3801 38335
rect 3801 38301 3835 38335
rect 3835 38301 3844 38335
rect 3792 38292 3844 38301
rect 4896 38292 4948 38344
rect 6368 38292 6420 38344
rect 9680 38335 9732 38344
rect 9680 38301 9689 38335
rect 9689 38301 9723 38335
rect 9723 38301 9732 38335
rect 9680 38292 9732 38301
rect 10232 38292 10284 38344
rect 11796 38360 11848 38412
rect 13820 38360 13872 38412
rect 11612 38335 11664 38344
rect 11612 38301 11621 38335
rect 11621 38301 11655 38335
rect 11655 38301 11664 38335
rect 11612 38292 11664 38301
rect 12256 38292 12308 38344
rect 12532 38292 12584 38344
rect 13360 38335 13412 38344
rect 13360 38301 13369 38335
rect 13369 38301 13403 38335
rect 13403 38301 13412 38335
rect 13360 38292 13412 38301
rect 5540 38267 5592 38276
rect 5540 38233 5574 38267
rect 5574 38233 5592 38267
rect 5540 38224 5592 38233
rect 5632 38224 5684 38276
rect 4252 38156 4304 38208
rect 10600 38156 10652 38208
rect 12256 38156 12308 38208
rect 6880 38054 6932 38106
rect 6944 38054 6996 38106
rect 7008 38054 7060 38106
rect 7072 38054 7124 38106
rect 7136 38054 7188 38106
rect 12811 38054 12863 38106
rect 12875 38054 12927 38106
rect 12939 38054 12991 38106
rect 13003 38054 13055 38106
rect 13067 38054 13119 38106
rect 8208 37952 8260 38004
rect 9680 37952 9732 38004
rect 12532 37952 12584 38004
rect 2780 37816 2832 37868
rect 5632 37884 5684 37936
rect 6736 37884 6788 37936
rect 4712 37816 4764 37868
rect 6552 37816 6604 37868
rect 8760 37884 8812 37936
rect 10692 37884 10744 37936
rect 10876 37884 10928 37936
rect 3148 37791 3200 37800
rect 3148 37757 3157 37791
rect 3157 37757 3191 37791
rect 3191 37757 3200 37791
rect 3148 37748 3200 37757
rect 7380 37816 7432 37868
rect 7748 37816 7800 37868
rect 8852 37859 8904 37868
rect 8852 37825 8861 37859
rect 8861 37825 8895 37859
rect 8895 37825 8904 37859
rect 8852 37816 8904 37825
rect 8024 37748 8076 37800
rect 8300 37748 8352 37800
rect 9772 37859 9824 37868
rect 9772 37825 9786 37859
rect 9786 37825 9820 37859
rect 9820 37825 9824 37859
rect 9772 37816 9824 37825
rect 10600 37859 10652 37868
rect 10232 37748 10284 37800
rect 10600 37825 10609 37859
rect 10609 37825 10643 37859
rect 10643 37825 10652 37859
rect 10600 37816 10652 37825
rect 13820 37884 13872 37936
rect 11796 37859 11848 37868
rect 11796 37825 11830 37859
rect 11830 37825 11848 37859
rect 14004 37859 14056 37868
rect 11796 37816 11848 37825
rect 14004 37825 14013 37859
rect 14013 37825 14047 37859
rect 14047 37825 14056 37859
rect 14004 37816 14056 37825
rect 14188 37859 14240 37868
rect 14188 37825 14197 37859
rect 14197 37825 14231 37859
rect 14231 37825 14240 37859
rect 14188 37816 14240 37825
rect 10692 37748 10744 37800
rect 10968 37748 11020 37800
rect 13360 37748 13412 37800
rect 2964 37655 3016 37664
rect 2964 37621 2973 37655
rect 2973 37621 3007 37655
rect 3007 37621 3016 37655
rect 2964 37612 3016 37621
rect 5080 37612 5132 37664
rect 5356 37612 5408 37664
rect 9404 37612 9456 37664
rect 10416 37655 10468 37664
rect 10416 37621 10425 37655
rect 10425 37621 10459 37655
rect 10459 37621 10468 37655
rect 10416 37612 10468 37621
rect 3915 37510 3967 37562
rect 3979 37510 4031 37562
rect 4043 37510 4095 37562
rect 4107 37510 4159 37562
rect 4171 37510 4223 37562
rect 9846 37510 9898 37562
rect 9910 37510 9962 37562
rect 9974 37510 10026 37562
rect 10038 37510 10090 37562
rect 10102 37510 10154 37562
rect 15776 37510 15828 37562
rect 15840 37510 15892 37562
rect 15904 37510 15956 37562
rect 15968 37510 16020 37562
rect 16032 37510 16084 37562
rect 6644 37451 6696 37460
rect 6644 37417 6653 37451
rect 6653 37417 6687 37451
rect 6687 37417 6696 37451
rect 6644 37408 6696 37417
rect 7288 37408 7340 37460
rect 10416 37451 10468 37460
rect 10416 37417 10425 37451
rect 10425 37417 10459 37451
rect 10459 37417 10468 37451
rect 10416 37408 10468 37417
rect 11796 37451 11848 37460
rect 11796 37417 11805 37451
rect 11805 37417 11839 37451
rect 11839 37417 11848 37451
rect 11796 37408 11848 37417
rect 3148 37204 3200 37256
rect 4896 37340 4948 37392
rect 7564 37340 7616 37392
rect 7932 37340 7984 37392
rect 8208 37340 8260 37392
rect 9772 37340 9824 37392
rect 4988 37315 5040 37324
rect 4988 37281 4997 37315
rect 4997 37281 5031 37315
rect 5031 37281 5040 37315
rect 4988 37272 5040 37281
rect 7472 37272 7524 37324
rect 10876 37340 10928 37392
rect 10692 37272 10744 37324
rect 2780 37068 2832 37120
rect 3608 37136 3660 37188
rect 3700 37136 3752 37188
rect 4252 37247 4304 37256
rect 4252 37213 4261 37247
rect 4261 37213 4295 37247
rect 4295 37213 4304 37247
rect 4252 37204 4304 37213
rect 4436 37247 4488 37256
rect 4436 37213 4445 37247
rect 4445 37213 4479 37247
rect 4479 37213 4488 37247
rect 5080 37247 5132 37256
rect 4436 37204 4488 37213
rect 5080 37213 5089 37247
rect 5089 37213 5123 37247
rect 5123 37213 5132 37247
rect 5080 37204 5132 37213
rect 4528 37136 4580 37188
rect 5540 37136 5592 37188
rect 5724 37136 5776 37188
rect 6460 37136 6512 37188
rect 9128 37204 9180 37256
rect 10508 37247 10560 37256
rect 7288 37179 7340 37188
rect 7288 37145 7297 37179
rect 7297 37145 7331 37179
rect 7331 37145 7340 37179
rect 7288 37136 7340 37145
rect 7564 37136 7616 37188
rect 7840 37179 7892 37188
rect 7840 37145 7849 37179
rect 7849 37145 7883 37179
rect 7883 37145 7892 37179
rect 7840 37136 7892 37145
rect 8300 37136 8352 37188
rect 10508 37213 10517 37247
rect 10517 37213 10551 37247
rect 10551 37213 10560 37247
rect 10508 37204 10560 37213
rect 11152 37247 11204 37256
rect 11152 37213 11161 37247
rect 11161 37213 11195 37247
rect 11195 37213 11204 37247
rect 11152 37204 11204 37213
rect 12256 37247 12308 37256
rect 5448 37111 5500 37120
rect 5448 37077 5457 37111
rect 5457 37077 5491 37111
rect 5491 37077 5500 37111
rect 5448 37068 5500 37077
rect 7932 37111 7984 37120
rect 7932 37077 7947 37111
rect 7947 37077 7981 37111
rect 7981 37077 7984 37111
rect 7932 37068 7984 37077
rect 12256 37213 12265 37247
rect 12265 37213 12299 37247
rect 12299 37213 12308 37247
rect 12256 37204 12308 37213
rect 12532 37136 12584 37188
rect 12348 37068 12400 37120
rect 13268 37204 13320 37256
rect 6880 36966 6932 37018
rect 6944 36966 6996 37018
rect 7008 36966 7060 37018
rect 7072 36966 7124 37018
rect 7136 36966 7188 37018
rect 12811 36966 12863 37018
rect 12875 36966 12927 37018
rect 12939 36966 12991 37018
rect 13003 36966 13055 37018
rect 13067 36966 13119 37018
rect 3792 36864 3844 36916
rect 4988 36864 5040 36916
rect 6552 36907 6604 36916
rect 6552 36873 6561 36907
rect 6561 36873 6595 36907
rect 6595 36873 6604 36907
rect 6552 36864 6604 36873
rect 4712 36839 4764 36848
rect 4712 36805 4721 36839
rect 4721 36805 4755 36839
rect 4755 36805 4764 36839
rect 4712 36796 4764 36805
rect 5448 36796 5500 36848
rect 2780 36728 2832 36780
rect 2688 36660 2740 36712
rect 2964 36660 3016 36712
rect 3608 36660 3660 36712
rect 4620 36660 4672 36712
rect 5080 36771 5132 36780
rect 5080 36737 5089 36771
rect 5089 36737 5123 36771
rect 5123 36737 5132 36771
rect 5080 36728 5132 36737
rect 5356 36728 5408 36780
rect 7472 36864 7524 36916
rect 10232 36864 10284 36916
rect 13820 36864 13872 36916
rect 7380 36796 7432 36848
rect 8116 36796 8168 36848
rect 7840 36728 7892 36780
rect 9404 36771 9456 36780
rect 9404 36737 9438 36771
rect 9438 36737 9456 36771
rect 9404 36728 9456 36737
rect 12716 36728 12768 36780
rect 15384 36728 15436 36780
rect 15568 36771 15620 36780
rect 15568 36737 15577 36771
rect 15577 36737 15611 36771
rect 15611 36737 15620 36771
rect 15568 36728 15620 36737
rect 16580 36660 16632 36712
rect 17408 36660 17460 36712
rect 5632 36592 5684 36644
rect 4896 36567 4948 36576
rect 4896 36533 4905 36567
rect 4905 36533 4939 36567
rect 4939 36533 4948 36567
rect 4896 36524 4948 36533
rect 15384 36567 15436 36576
rect 15384 36533 15393 36567
rect 15393 36533 15427 36567
rect 15427 36533 15436 36567
rect 15384 36524 15436 36533
rect 3915 36422 3967 36474
rect 3979 36422 4031 36474
rect 4043 36422 4095 36474
rect 4107 36422 4159 36474
rect 4171 36422 4223 36474
rect 9846 36422 9898 36474
rect 9910 36422 9962 36474
rect 9974 36422 10026 36474
rect 10038 36422 10090 36474
rect 10102 36422 10154 36474
rect 15776 36422 15828 36474
rect 15840 36422 15892 36474
rect 15904 36422 15956 36474
rect 15968 36422 16020 36474
rect 16032 36422 16084 36474
rect 3148 36320 3200 36372
rect 4896 36320 4948 36372
rect 7840 36363 7892 36372
rect 7840 36329 7849 36363
rect 7849 36329 7883 36363
rect 7883 36329 7892 36363
rect 7840 36320 7892 36329
rect 10508 36320 10560 36372
rect 8392 36252 8444 36304
rect 16580 36252 16632 36304
rect 4528 36184 4580 36236
rect 8116 36184 8168 36236
rect 3608 36048 3660 36100
rect 5356 36116 5408 36168
rect 7932 36116 7984 36168
rect 8300 36159 8352 36168
rect 8300 36125 8309 36159
rect 8309 36125 8343 36159
rect 8343 36125 8352 36159
rect 8300 36116 8352 36125
rect 10600 36116 10652 36168
rect 10968 36159 11020 36168
rect 10968 36125 10977 36159
rect 10977 36125 11011 36159
rect 11011 36125 11020 36159
rect 10968 36116 11020 36125
rect 14924 36159 14976 36168
rect 14924 36125 14933 36159
rect 14933 36125 14967 36159
rect 14967 36125 14976 36159
rect 14924 36116 14976 36125
rect 16488 36116 16540 36168
rect 4804 36048 4856 36100
rect 9220 36091 9272 36100
rect 9220 36057 9254 36091
rect 9254 36057 9272 36091
rect 9220 36048 9272 36057
rect 8852 35980 8904 36032
rect 14740 36023 14792 36032
rect 14740 35989 14749 36023
rect 14749 35989 14783 36023
rect 14783 35989 14792 36023
rect 14740 35980 14792 35989
rect 15200 35980 15252 36032
rect 15660 35980 15712 36032
rect 16120 35980 16172 36032
rect 16764 35980 16816 36032
rect 6880 35878 6932 35930
rect 6944 35878 6996 35930
rect 7008 35878 7060 35930
rect 7072 35878 7124 35930
rect 7136 35878 7188 35930
rect 12811 35878 12863 35930
rect 12875 35878 12927 35930
rect 12939 35878 12991 35930
rect 13003 35878 13055 35930
rect 13067 35878 13119 35930
rect 9220 35776 9272 35828
rect 16488 35776 16540 35828
rect 4528 35640 4580 35692
rect 8852 35640 8904 35692
rect 9404 35683 9456 35692
rect 9404 35649 9413 35683
rect 9413 35649 9447 35683
rect 9447 35649 9456 35683
rect 9404 35640 9456 35649
rect 1400 35615 1452 35624
rect 1400 35581 1409 35615
rect 1409 35581 1443 35615
rect 1443 35581 1452 35615
rect 1400 35572 1452 35581
rect 1676 35615 1728 35624
rect 1676 35581 1685 35615
rect 1685 35581 1719 35615
rect 1719 35581 1728 35615
rect 1676 35572 1728 35581
rect 8392 35572 8444 35624
rect 9588 35683 9640 35692
rect 9588 35649 9597 35683
rect 9597 35649 9631 35683
rect 9631 35649 9640 35683
rect 9588 35640 9640 35649
rect 10600 35640 10652 35692
rect 11152 35640 11204 35692
rect 15384 35640 15436 35692
rect 9680 35572 9732 35624
rect 13820 35572 13872 35624
rect 14556 35572 14608 35624
rect 5724 35436 5776 35488
rect 15660 35436 15712 35488
rect 17408 35640 17460 35692
rect 16764 35615 16816 35624
rect 16764 35581 16773 35615
rect 16773 35581 16807 35615
rect 16807 35581 16816 35615
rect 16764 35572 16816 35581
rect 16304 35436 16356 35488
rect 3915 35334 3967 35386
rect 3979 35334 4031 35386
rect 4043 35334 4095 35386
rect 4107 35334 4159 35386
rect 4171 35334 4223 35386
rect 9846 35334 9898 35386
rect 9910 35334 9962 35386
rect 9974 35334 10026 35386
rect 10038 35334 10090 35386
rect 10102 35334 10154 35386
rect 15776 35334 15828 35386
rect 15840 35334 15892 35386
rect 15904 35334 15956 35386
rect 15968 35334 16020 35386
rect 16032 35334 16084 35386
rect 16764 35275 16816 35284
rect 16764 35241 16773 35275
rect 16773 35241 16807 35275
rect 16807 35241 16816 35275
rect 16764 35232 16816 35241
rect 7288 35164 7340 35216
rect 14372 35071 14424 35080
rect 14372 35037 14381 35071
rect 14381 35037 14415 35071
rect 14415 35037 14424 35071
rect 14372 35028 14424 35037
rect 15200 35164 15252 35216
rect 14556 35096 14608 35148
rect 14740 35028 14792 35080
rect 14832 35071 14884 35080
rect 14832 35037 14841 35071
rect 14841 35037 14875 35071
rect 14875 35037 14884 35071
rect 14832 35028 14884 35037
rect 10416 34960 10468 35012
rect 14188 34935 14240 34944
rect 14188 34901 14197 34935
rect 14197 34901 14231 34935
rect 14231 34901 14240 34935
rect 14188 34892 14240 34901
rect 16672 34960 16724 35012
rect 16304 34892 16356 34944
rect 6880 34790 6932 34842
rect 6944 34790 6996 34842
rect 7008 34790 7060 34842
rect 7072 34790 7124 34842
rect 7136 34790 7188 34842
rect 12811 34790 12863 34842
rect 12875 34790 12927 34842
rect 12939 34790 12991 34842
rect 13003 34790 13055 34842
rect 13067 34790 13119 34842
rect 10416 34731 10468 34740
rect 10416 34697 10425 34731
rect 10425 34697 10459 34731
rect 10459 34697 10468 34731
rect 16672 34731 16724 34740
rect 10416 34688 10468 34697
rect 16672 34697 16681 34731
rect 16681 34697 16715 34731
rect 16715 34697 16724 34731
rect 16672 34688 16724 34697
rect 14188 34620 14240 34672
rect 10508 34595 10560 34604
rect 10508 34561 10517 34595
rect 10517 34561 10551 34595
rect 10551 34561 10560 34595
rect 10508 34552 10560 34561
rect 11796 34595 11848 34604
rect 11796 34561 11805 34595
rect 11805 34561 11839 34595
rect 11839 34561 11848 34595
rect 11796 34552 11848 34561
rect 14556 34595 14608 34604
rect 11520 34484 11572 34536
rect 14556 34561 14565 34595
rect 14565 34561 14599 34595
rect 14599 34561 14608 34595
rect 14556 34552 14608 34561
rect 15568 34552 15620 34604
rect 16856 34595 16908 34604
rect 16856 34561 16865 34595
rect 16865 34561 16899 34595
rect 16899 34561 16908 34595
rect 16856 34552 16908 34561
rect 12716 34527 12768 34536
rect 12716 34493 12725 34527
rect 12725 34493 12759 34527
rect 12759 34493 12768 34527
rect 12716 34484 12768 34493
rect 15016 34527 15068 34536
rect 15016 34493 15025 34527
rect 15025 34493 15059 34527
rect 15059 34493 15068 34527
rect 15016 34484 15068 34493
rect 11980 34391 12032 34400
rect 11980 34357 11989 34391
rect 11989 34357 12023 34391
rect 12023 34357 12032 34391
rect 11980 34348 12032 34357
rect 13176 34391 13228 34400
rect 13176 34357 13185 34391
rect 13185 34357 13219 34391
rect 13219 34357 13228 34391
rect 13176 34348 13228 34357
rect 3915 34246 3967 34298
rect 3979 34246 4031 34298
rect 4043 34246 4095 34298
rect 4107 34246 4159 34298
rect 4171 34246 4223 34298
rect 9846 34246 9898 34298
rect 9910 34246 9962 34298
rect 9974 34246 10026 34298
rect 10038 34246 10090 34298
rect 10102 34246 10154 34298
rect 15776 34246 15828 34298
rect 15840 34246 15892 34298
rect 15904 34246 15956 34298
rect 15968 34246 16020 34298
rect 16032 34246 16084 34298
rect 8024 34144 8076 34196
rect 5908 33940 5960 33992
rect 6460 33940 6512 33992
rect 7564 33940 7616 33992
rect 9128 33940 9180 33992
rect 13360 33983 13412 33992
rect 13360 33949 13369 33983
rect 13369 33949 13403 33983
rect 13403 33949 13412 33983
rect 13360 33940 13412 33949
rect 14096 33983 14148 33992
rect 14096 33949 14105 33983
rect 14105 33949 14139 33983
rect 14139 33949 14148 33983
rect 14096 33940 14148 33949
rect 7472 33872 7524 33924
rect 8024 33872 8076 33924
rect 14832 34144 14884 34196
rect 16856 34144 16908 34196
rect 15660 34051 15712 34060
rect 15660 34017 15669 34051
rect 15669 34017 15703 34051
rect 15703 34017 15712 34051
rect 15660 34008 15712 34017
rect 15384 33872 15436 33924
rect 5908 33847 5960 33856
rect 5908 33813 5923 33847
rect 5923 33813 5957 33847
rect 5957 33813 5960 33847
rect 5908 33804 5960 33813
rect 6644 33847 6696 33856
rect 6644 33813 6653 33847
rect 6653 33813 6687 33847
rect 6687 33813 6696 33847
rect 6644 33804 6696 33813
rect 11796 33804 11848 33856
rect 6880 33702 6932 33754
rect 6944 33702 6996 33754
rect 7008 33702 7060 33754
rect 7072 33702 7124 33754
rect 7136 33702 7188 33754
rect 12811 33702 12863 33754
rect 12875 33702 12927 33754
rect 12939 33702 12991 33754
rect 13003 33702 13055 33754
rect 13067 33702 13119 33754
rect 5908 33532 5960 33584
rect 7288 33532 7340 33584
rect 8300 33532 8352 33584
rect 8116 33507 8168 33516
rect 8116 33473 8125 33507
rect 8125 33473 8159 33507
rect 8159 33473 8168 33507
rect 8116 33464 8168 33473
rect 8208 33507 8260 33516
rect 8208 33473 8217 33507
rect 8217 33473 8251 33507
rect 8251 33473 8260 33507
rect 11796 33532 11848 33584
rect 13176 33575 13228 33584
rect 13176 33541 13185 33575
rect 13185 33541 13219 33575
rect 13219 33541 13228 33575
rect 13176 33532 13228 33541
rect 8208 33464 8260 33473
rect 5816 33396 5868 33448
rect 11520 33464 11572 33516
rect 7380 33371 7432 33380
rect 4436 33260 4488 33312
rect 7380 33337 7389 33371
rect 7389 33337 7423 33371
rect 7423 33337 7432 33371
rect 7380 33328 7432 33337
rect 9220 33396 9272 33448
rect 10416 33396 10468 33448
rect 11980 33507 12032 33516
rect 11980 33473 11989 33507
rect 11989 33473 12023 33507
rect 12023 33473 12032 33507
rect 11980 33464 12032 33473
rect 12256 33507 12308 33516
rect 12256 33473 12265 33507
rect 12265 33473 12299 33507
rect 12299 33473 12308 33507
rect 12256 33464 12308 33473
rect 14004 33464 14056 33516
rect 14372 33464 14424 33516
rect 12072 33396 12124 33448
rect 15016 33439 15068 33448
rect 15016 33405 15025 33439
rect 15025 33405 15059 33439
rect 15059 33405 15068 33439
rect 15016 33396 15068 33405
rect 8760 33328 8812 33380
rect 12440 33328 12492 33380
rect 5816 33303 5868 33312
rect 5816 33269 5825 33303
rect 5825 33269 5859 33303
rect 5859 33269 5868 33303
rect 5816 33260 5868 33269
rect 6460 33260 6512 33312
rect 8944 33303 8996 33312
rect 8944 33269 8953 33303
rect 8953 33269 8987 33303
rect 8987 33269 8996 33303
rect 8944 33260 8996 33269
rect 10232 33260 10284 33312
rect 11888 33260 11940 33312
rect 3915 33158 3967 33210
rect 3979 33158 4031 33210
rect 4043 33158 4095 33210
rect 4107 33158 4159 33210
rect 4171 33158 4223 33210
rect 9846 33158 9898 33210
rect 9910 33158 9962 33210
rect 9974 33158 10026 33210
rect 10038 33158 10090 33210
rect 10102 33158 10154 33210
rect 15776 33158 15828 33210
rect 15840 33158 15892 33210
rect 15904 33158 15956 33210
rect 15968 33158 16020 33210
rect 16032 33158 16084 33210
rect 4712 33056 4764 33108
rect 3700 32852 3752 32904
rect 5080 32988 5132 33040
rect 8300 33056 8352 33108
rect 8944 33056 8996 33108
rect 10692 33056 10744 33108
rect 11520 33099 11572 33108
rect 11520 33065 11529 33099
rect 11529 33065 11563 33099
rect 11563 33065 11572 33099
rect 11520 33056 11572 33065
rect 14096 33099 14148 33108
rect 14096 33065 14105 33099
rect 14105 33065 14139 33099
rect 14139 33065 14148 33099
rect 14096 33056 14148 33065
rect 9680 32988 9732 33040
rect 10416 32988 10468 33040
rect 4620 32920 4672 32972
rect 4528 32852 4580 32904
rect 4712 32895 4764 32904
rect 4712 32861 4721 32895
rect 4721 32861 4755 32895
rect 4755 32861 4764 32895
rect 4712 32852 4764 32861
rect 4252 32827 4304 32836
rect 3884 32716 3936 32768
rect 4252 32793 4261 32827
rect 4261 32793 4295 32827
rect 4295 32793 4304 32827
rect 4252 32784 4304 32793
rect 5080 32852 5132 32904
rect 5632 32920 5684 32972
rect 8208 32920 8260 32972
rect 9036 32920 9088 32972
rect 5816 32852 5868 32904
rect 7380 32852 7432 32904
rect 6644 32784 6696 32836
rect 8392 32852 8444 32904
rect 9128 32895 9180 32904
rect 9128 32861 9137 32895
rect 9137 32861 9171 32895
rect 9171 32861 9180 32895
rect 9128 32852 9180 32861
rect 10232 32920 10284 32972
rect 13176 32920 13228 32972
rect 15384 32963 15436 32972
rect 15384 32929 15393 32963
rect 15393 32929 15427 32963
rect 15427 32929 15436 32963
rect 15384 32920 15436 32929
rect 16764 32920 16816 32972
rect 13360 32852 13412 32904
rect 13728 32852 13780 32904
rect 14188 32852 14240 32904
rect 15016 32852 15068 32904
rect 8116 32784 8168 32836
rect 10784 32784 10836 32836
rect 12624 32827 12676 32836
rect 12624 32793 12642 32827
rect 12642 32793 12676 32827
rect 12624 32784 12676 32793
rect 4620 32716 4672 32768
rect 6184 32716 6236 32768
rect 7288 32716 7340 32768
rect 6880 32614 6932 32666
rect 6944 32614 6996 32666
rect 7008 32614 7060 32666
rect 7072 32614 7124 32666
rect 7136 32614 7188 32666
rect 12811 32614 12863 32666
rect 12875 32614 12927 32666
rect 12939 32614 12991 32666
rect 13003 32614 13055 32666
rect 13067 32614 13119 32666
rect 6460 32555 6512 32564
rect 6460 32521 6469 32555
rect 6469 32521 6503 32555
rect 6503 32521 6512 32555
rect 6460 32512 6512 32521
rect 7564 32555 7616 32564
rect 4436 32444 4488 32496
rect 3884 32419 3936 32428
rect 3884 32385 3918 32419
rect 3918 32385 3936 32419
rect 3884 32376 3936 32385
rect 6000 32444 6052 32496
rect 6092 32444 6144 32496
rect 7104 32444 7156 32496
rect 7564 32521 7573 32555
rect 7573 32521 7607 32555
rect 7607 32521 7616 32555
rect 7564 32512 7616 32521
rect 8852 32555 8904 32564
rect 8852 32521 8861 32555
rect 8861 32521 8895 32555
rect 8895 32521 8904 32555
rect 8852 32512 8904 32521
rect 10324 32512 10376 32564
rect 11888 32512 11940 32564
rect 7932 32444 7984 32496
rect 8392 32444 8444 32496
rect 7288 32419 7340 32428
rect 7288 32385 7298 32419
rect 7298 32385 7332 32419
rect 7332 32385 7340 32419
rect 7288 32376 7340 32385
rect 8116 32376 8168 32428
rect 9680 32444 9732 32496
rect 10232 32444 10284 32496
rect 10784 32487 10836 32496
rect 10784 32453 10793 32487
rect 10793 32453 10827 32487
rect 10827 32453 10836 32487
rect 10784 32444 10836 32453
rect 12716 32444 12768 32496
rect 7472 32308 7524 32360
rect 8208 32308 8260 32360
rect 8392 32308 8444 32360
rect 11888 32419 11940 32428
rect 11888 32385 11897 32419
rect 11897 32385 11931 32419
rect 11931 32385 11940 32419
rect 11888 32376 11940 32385
rect 12072 32376 12124 32428
rect 12256 32419 12308 32428
rect 12256 32385 12265 32419
rect 12265 32385 12299 32419
rect 12299 32385 12308 32419
rect 12256 32376 12308 32385
rect 12440 32308 12492 32360
rect 7288 32240 7340 32292
rect 11980 32240 12032 32292
rect 13176 32240 13228 32292
rect 4988 32215 5040 32224
rect 4988 32181 4997 32215
rect 4997 32181 5031 32215
rect 5031 32181 5040 32215
rect 4988 32172 5040 32181
rect 6920 32172 6972 32224
rect 10876 32215 10928 32224
rect 10876 32181 10885 32215
rect 10885 32181 10919 32215
rect 10919 32181 10928 32215
rect 10876 32172 10928 32181
rect 12348 32172 12400 32224
rect 13728 32172 13780 32224
rect 3915 32070 3967 32122
rect 3979 32070 4031 32122
rect 4043 32070 4095 32122
rect 4107 32070 4159 32122
rect 4171 32070 4223 32122
rect 9846 32070 9898 32122
rect 9910 32070 9962 32122
rect 9974 32070 10026 32122
rect 10038 32070 10090 32122
rect 10102 32070 10154 32122
rect 15776 32070 15828 32122
rect 15840 32070 15892 32122
rect 15904 32070 15956 32122
rect 15968 32070 16020 32122
rect 16032 32070 16084 32122
rect 4252 32011 4304 32020
rect 4252 31977 4261 32011
rect 4261 31977 4295 32011
rect 4295 31977 4304 32011
rect 4252 31968 4304 31977
rect 4528 31968 4580 32020
rect 5080 31968 5132 32020
rect 7472 31968 7524 32020
rect 9588 31968 9640 32020
rect 12624 31968 12676 32020
rect 3792 31832 3844 31884
rect 5816 31875 5868 31884
rect 5816 31841 5825 31875
rect 5825 31841 5859 31875
rect 5859 31841 5868 31875
rect 5816 31832 5868 31841
rect 7012 31900 7064 31952
rect 3976 31807 4028 31816
rect 3976 31773 3985 31807
rect 3985 31773 4019 31807
rect 4019 31773 4028 31807
rect 3976 31764 4028 31773
rect 4804 31807 4856 31816
rect 4804 31773 4813 31807
rect 4813 31773 4847 31807
rect 4847 31773 4856 31807
rect 4804 31764 4856 31773
rect 4988 31807 5040 31816
rect 4988 31773 4997 31807
rect 4997 31773 5031 31807
rect 5031 31773 5040 31807
rect 5632 31807 5684 31816
rect 4988 31764 5040 31773
rect 5632 31773 5641 31807
rect 5641 31773 5675 31807
rect 5675 31773 5684 31807
rect 5632 31764 5684 31773
rect 5724 31764 5776 31816
rect 6092 31764 6144 31816
rect 9404 31832 9456 31884
rect 5448 31696 5500 31748
rect 6736 31807 6788 31816
rect 6736 31773 6746 31807
rect 6746 31773 6780 31807
rect 6780 31773 6788 31807
rect 7012 31807 7064 31816
rect 6736 31764 6788 31773
rect 7012 31773 7021 31807
rect 7021 31773 7055 31807
rect 7055 31773 7064 31807
rect 7012 31764 7064 31773
rect 7104 31807 7156 31816
rect 7104 31773 7118 31807
rect 7118 31773 7152 31807
rect 7152 31773 7156 31807
rect 7932 31807 7984 31816
rect 7104 31764 7156 31773
rect 7932 31773 7941 31807
rect 7941 31773 7975 31807
rect 7975 31773 7984 31807
rect 7932 31764 7984 31773
rect 10324 31832 10376 31884
rect 10416 31832 10468 31884
rect 10784 31832 10836 31884
rect 12440 31832 12492 31884
rect 6920 31739 6972 31748
rect 6920 31705 6929 31739
rect 6929 31705 6963 31739
rect 6963 31705 6972 31739
rect 6920 31696 6972 31705
rect 7840 31628 7892 31680
rect 10416 31696 10468 31748
rect 11796 31764 11848 31816
rect 11152 31696 11204 31748
rect 9956 31628 10008 31680
rect 6880 31526 6932 31578
rect 6944 31526 6996 31578
rect 7008 31526 7060 31578
rect 7072 31526 7124 31578
rect 7136 31526 7188 31578
rect 12811 31526 12863 31578
rect 12875 31526 12927 31578
rect 12939 31526 12991 31578
rect 13003 31526 13055 31578
rect 13067 31526 13119 31578
rect 3056 31424 3108 31476
rect 3976 31424 4028 31476
rect 5632 31424 5684 31476
rect 6736 31424 6788 31476
rect 4988 31288 5040 31340
rect 7288 31356 7340 31408
rect 9128 31356 9180 31408
rect 2596 31263 2648 31272
rect 2596 31229 2605 31263
rect 2605 31229 2639 31263
rect 2639 31229 2648 31263
rect 2596 31220 2648 31229
rect 3608 31220 3660 31272
rect 7840 31220 7892 31272
rect 8760 31331 8812 31340
rect 8760 31297 8769 31331
rect 8769 31297 8803 31331
rect 8803 31297 8812 31331
rect 8760 31288 8812 31297
rect 10140 31424 10192 31476
rect 10968 31424 11020 31476
rect 9956 31331 10008 31340
rect 9956 31297 9965 31331
rect 9965 31297 9999 31331
rect 9999 31297 10008 31331
rect 9956 31288 10008 31297
rect 8852 31220 8904 31272
rect 9588 31220 9640 31272
rect 10324 31288 10376 31340
rect 10600 31288 10652 31340
rect 11152 31288 11204 31340
rect 14188 31288 14240 31340
rect 14372 31331 14424 31340
rect 14372 31297 14381 31331
rect 14381 31297 14415 31331
rect 14415 31297 14424 31331
rect 14372 31288 14424 31297
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 10232 31220 10284 31272
rect 14280 31220 14332 31272
rect 9772 31152 9824 31204
rect 10600 31152 10652 31204
rect 3516 31084 3568 31136
rect 4252 31127 4304 31136
rect 4252 31093 4261 31127
rect 4261 31093 4295 31127
rect 4295 31093 4304 31127
rect 6828 31127 6880 31136
rect 4252 31084 4304 31093
rect 6828 31093 6837 31127
rect 6837 31093 6871 31127
rect 6871 31093 6880 31127
rect 6828 31084 6880 31093
rect 7196 31127 7248 31136
rect 7196 31093 7205 31127
rect 7205 31093 7239 31127
rect 7239 31093 7248 31127
rect 7196 31084 7248 31093
rect 7932 31084 7984 31136
rect 8300 31127 8352 31136
rect 8300 31093 8309 31127
rect 8309 31093 8343 31127
rect 8343 31093 8352 31127
rect 8300 31084 8352 31093
rect 10968 31084 11020 31136
rect 13360 31084 13412 31136
rect 16672 31127 16724 31136
rect 16672 31093 16681 31127
rect 16681 31093 16715 31127
rect 16715 31093 16724 31127
rect 16672 31084 16724 31093
rect 3915 30982 3967 31034
rect 3979 30982 4031 31034
rect 4043 30982 4095 31034
rect 4107 30982 4159 31034
rect 4171 30982 4223 31034
rect 9846 30982 9898 31034
rect 9910 30982 9962 31034
rect 9974 30982 10026 31034
rect 10038 30982 10090 31034
rect 10102 30982 10154 31034
rect 15776 30982 15828 31034
rect 15840 30982 15892 31034
rect 15904 30982 15956 31034
rect 15968 30982 16020 31034
rect 16032 30982 16084 31034
rect 2688 30923 2740 30932
rect 2688 30889 2697 30923
rect 2697 30889 2731 30923
rect 2731 30889 2740 30923
rect 2688 30880 2740 30889
rect 3792 30880 3844 30932
rect 8392 30880 8444 30932
rect 10416 30880 10468 30932
rect 3056 30855 3108 30864
rect 3056 30821 3065 30855
rect 3065 30821 3099 30855
rect 3099 30821 3108 30855
rect 3056 30812 3108 30821
rect 10784 30787 10836 30796
rect 10784 30753 10793 30787
rect 10793 30753 10827 30787
rect 10827 30753 10836 30787
rect 10784 30744 10836 30753
rect 2872 30719 2924 30728
rect 2872 30685 2881 30719
rect 2881 30685 2915 30719
rect 2915 30685 2924 30719
rect 2872 30676 2924 30685
rect 2964 30719 3016 30728
rect 2964 30685 2973 30719
rect 2973 30685 3007 30719
rect 3007 30685 3016 30719
rect 2964 30676 3016 30685
rect 3516 30676 3568 30728
rect 3608 30676 3660 30728
rect 7288 30676 7340 30728
rect 9036 30676 9088 30728
rect 6828 30608 6880 30660
rect 7196 30608 7248 30660
rect 7380 30608 7432 30660
rect 7748 30608 7800 30660
rect 9588 30676 9640 30728
rect 10600 30719 10652 30728
rect 10600 30685 10609 30719
rect 10609 30685 10643 30719
rect 10643 30685 10652 30719
rect 13360 30719 13412 30728
rect 10600 30676 10652 30685
rect 13360 30685 13369 30719
rect 13369 30685 13403 30719
rect 13403 30685 13412 30719
rect 13360 30676 13412 30685
rect 15476 30719 15528 30728
rect 15476 30685 15485 30719
rect 15485 30685 15519 30719
rect 15519 30685 15528 30719
rect 15476 30676 15528 30685
rect 9680 30651 9732 30660
rect 3792 30540 3844 30592
rect 4252 30540 4304 30592
rect 7840 30583 7892 30592
rect 7840 30549 7849 30583
rect 7849 30549 7883 30583
rect 7883 30549 7892 30583
rect 7840 30540 7892 30549
rect 9680 30617 9689 30651
rect 9689 30617 9723 30651
rect 9723 30617 9732 30651
rect 9680 30608 9732 30617
rect 10968 30608 11020 30660
rect 15752 30608 15804 30660
rect 17500 30608 17552 30660
rect 9956 30540 10008 30592
rect 10416 30540 10468 30592
rect 14004 30540 14056 30592
rect 14280 30540 14332 30592
rect 16580 30540 16632 30592
rect 6880 30438 6932 30490
rect 6944 30438 6996 30490
rect 7008 30438 7060 30490
rect 7072 30438 7124 30490
rect 7136 30438 7188 30490
rect 12811 30438 12863 30490
rect 12875 30438 12927 30490
rect 12939 30438 12991 30490
rect 13003 30438 13055 30490
rect 13067 30438 13119 30490
rect 9036 30336 9088 30388
rect 15752 30379 15804 30388
rect 15752 30345 15761 30379
rect 15761 30345 15795 30379
rect 15795 30345 15804 30379
rect 15752 30336 15804 30345
rect 16856 30336 16908 30388
rect 17500 30379 17552 30388
rect 17500 30345 17509 30379
rect 17509 30345 17543 30379
rect 17543 30345 17552 30379
rect 17500 30336 17552 30345
rect 8300 30268 8352 30320
rect 9956 30268 10008 30320
rect 7288 30200 7340 30252
rect 9680 30200 9732 30252
rect 10232 30200 10284 30252
rect 10416 30200 10468 30252
rect 10784 30200 10836 30252
rect 11336 30132 11388 30184
rect 13728 30200 13780 30252
rect 15476 30268 15528 30320
rect 14004 30200 14056 30252
rect 14464 30200 14516 30252
rect 16764 30200 16816 30252
rect 16948 30200 17000 30252
rect 17684 30243 17736 30252
rect 17684 30209 17693 30243
rect 17693 30209 17727 30243
rect 17727 30209 17736 30243
rect 17684 30200 17736 30209
rect 16580 30132 16632 30184
rect 9680 29996 9732 30048
rect 10600 30039 10652 30048
rect 10600 30005 10609 30039
rect 10609 30005 10643 30039
rect 10643 30005 10652 30039
rect 10600 29996 10652 30005
rect 15108 29996 15160 30048
rect 3915 29894 3967 29946
rect 3979 29894 4031 29946
rect 4043 29894 4095 29946
rect 4107 29894 4159 29946
rect 4171 29894 4223 29946
rect 9846 29894 9898 29946
rect 9910 29894 9962 29946
rect 9974 29894 10026 29946
rect 10038 29894 10090 29946
rect 10102 29894 10154 29946
rect 15776 29894 15828 29946
rect 15840 29894 15892 29946
rect 15904 29894 15956 29946
rect 15968 29894 16020 29946
rect 16032 29894 16084 29946
rect 5448 29835 5500 29844
rect 5448 29801 5457 29835
rect 5457 29801 5491 29835
rect 5491 29801 5500 29835
rect 5448 29792 5500 29801
rect 12532 29792 12584 29844
rect 3792 29724 3844 29776
rect 2964 29656 3016 29708
rect 2872 29588 2924 29640
rect 7840 29656 7892 29708
rect 9680 29699 9732 29708
rect 9680 29665 9689 29699
rect 9689 29665 9723 29699
rect 9723 29665 9732 29699
rect 9680 29656 9732 29665
rect 13728 29792 13780 29844
rect 14464 29724 14516 29776
rect 14188 29656 14240 29708
rect 5632 29631 5684 29640
rect 5632 29597 5641 29631
rect 5641 29597 5675 29631
rect 5675 29597 5684 29631
rect 5632 29588 5684 29597
rect 5908 29631 5960 29640
rect 5908 29597 5917 29631
rect 5917 29597 5951 29631
rect 5951 29597 5960 29631
rect 5908 29588 5960 29597
rect 6092 29588 6144 29640
rect 6276 29588 6328 29640
rect 9588 29631 9640 29640
rect 9588 29597 9597 29631
rect 9597 29597 9631 29631
rect 9631 29597 9640 29631
rect 9588 29588 9640 29597
rect 10232 29588 10284 29640
rect 11336 29631 11388 29640
rect 11336 29597 11345 29631
rect 11345 29597 11379 29631
rect 11379 29597 11388 29631
rect 11336 29588 11388 29597
rect 13360 29631 13412 29640
rect 13360 29597 13369 29631
rect 13369 29597 13403 29631
rect 13403 29597 13412 29631
rect 13360 29588 13412 29597
rect 14280 29631 14332 29640
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 14372 29631 14424 29640
rect 14372 29597 14381 29631
rect 14381 29597 14415 29631
rect 14415 29597 14424 29631
rect 14372 29588 14424 29597
rect 9680 29520 9732 29572
rect 12072 29520 12124 29572
rect 14556 29563 14608 29572
rect 14556 29529 14565 29563
rect 14565 29529 14599 29563
rect 14599 29529 14608 29563
rect 15108 29588 15160 29640
rect 15476 29656 15528 29708
rect 14556 29520 14608 29529
rect 16672 29520 16724 29572
rect 10232 29452 10284 29504
rect 13636 29452 13688 29504
rect 15844 29452 15896 29504
rect 17592 29495 17644 29504
rect 17592 29461 17601 29495
rect 17601 29461 17635 29495
rect 17635 29461 17644 29495
rect 17592 29452 17644 29461
rect 6880 29350 6932 29402
rect 6944 29350 6996 29402
rect 7008 29350 7060 29402
rect 7072 29350 7124 29402
rect 7136 29350 7188 29402
rect 12811 29350 12863 29402
rect 12875 29350 12927 29402
rect 12939 29350 12991 29402
rect 13003 29350 13055 29402
rect 13067 29350 13119 29402
rect 2964 29248 3016 29300
rect 5908 29248 5960 29300
rect 14372 29248 14424 29300
rect 17684 29248 17736 29300
rect 2596 29087 2648 29096
rect 2596 29053 2605 29087
rect 2605 29053 2639 29087
rect 2639 29053 2648 29087
rect 2596 29044 2648 29053
rect 3792 29112 3844 29164
rect 2872 29044 2924 29096
rect 3332 29087 3384 29096
rect 3332 29053 3341 29087
rect 3341 29053 3375 29087
rect 3375 29053 3384 29087
rect 3332 29044 3384 29053
rect 4804 29044 4856 29096
rect 4160 28976 4212 29028
rect 15476 29112 15528 29164
rect 15844 29155 15896 29164
rect 15844 29121 15853 29155
rect 15853 29121 15887 29155
rect 15887 29121 15896 29155
rect 15844 29112 15896 29121
rect 16764 29155 16816 29164
rect 16764 29121 16773 29155
rect 16773 29121 16807 29155
rect 16807 29121 16816 29155
rect 16764 29112 16816 29121
rect 16948 29112 17000 29164
rect 5264 28976 5316 29028
rect 4252 28908 4304 28960
rect 3915 28806 3967 28858
rect 3979 28806 4031 28858
rect 4043 28806 4095 28858
rect 4107 28806 4159 28858
rect 4171 28806 4223 28858
rect 9846 28806 9898 28858
rect 9910 28806 9962 28858
rect 9974 28806 10026 28858
rect 10038 28806 10090 28858
rect 10102 28806 10154 28858
rect 15776 28806 15828 28858
rect 15840 28806 15892 28858
rect 15904 28806 15956 28858
rect 15968 28806 16020 28858
rect 16032 28806 16084 28858
rect 6276 28747 6328 28756
rect 6276 28713 6285 28747
rect 6285 28713 6319 28747
rect 6319 28713 6328 28747
rect 6276 28704 6328 28713
rect 12072 28747 12124 28756
rect 12072 28713 12081 28747
rect 12081 28713 12115 28747
rect 12115 28713 12124 28747
rect 12072 28704 12124 28713
rect 16764 28704 16816 28756
rect 14280 28636 14332 28688
rect 5908 28568 5960 28620
rect 3608 28500 3660 28552
rect 5540 28500 5592 28552
rect 12624 28568 12676 28620
rect 13728 28568 13780 28620
rect 6092 28543 6144 28552
rect 6092 28509 6101 28543
rect 6101 28509 6135 28543
rect 6135 28509 6144 28543
rect 6092 28500 6144 28509
rect 7380 28500 7432 28552
rect 7840 28500 7892 28552
rect 10232 28500 10284 28552
rect 10876 28500 10928 28552
rect 3792 28432 3844 28484
rect 5908 28475 5960 28484
rect 5908 28441 5917 28475
rect 5917 28441 5951 28475
rect 5951 28441 5960 28475
rect 5908 28432 5960 28441
rect 12348 28543 12400 28552
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 12716 28500 12768 28552
rect 13360 28500 13412 28552
rect 14372 28543 14424 28552
rect 14372 28509 14381 28543
rect 14381 28509 14415 28543
rect 14415 28509 14424 28543
rect 14372 28500 14424 28509
rect 15476 28568 15528 28620
rect 13544 28432 13596 28484
rect 13820 28432 13872 28484
rect 14556 28432 14608 28484
rect 16672 28432 16724 28484
rect 5264 28407 5316 28416
rect 5264 28373 5273 28407
rect 5273 28373 5307 28407
rect 5307 28373 5316 28407
rect 5264 28364 5316 28373
rect 7380 28407 7432 28416
rect 7380 28373 7389 28407
rect 7389 28373 7423 28407
rect 7423 28373 7432 28407
rect 7380 28364 7432 28373
rect 10232 28407 10284 28416
rect 10232 28373 10241 28407
rect 10241 28373 10275 28407
rect 10275 28373 10284 28407
rect 10232 28364 10284 28373
rect 14004 28364 14056 28416
rect 6880 28262 6932 28314
rect 6944 28262 6996 28314
rect 7008 28262 7060 28314
rect 7072 28262 7124 28314
rect 7136 28262 7188 28314
rect 12811 28262 12863 28314
rect 12875 28262 12927 28314
rect 12939 28262 12991 28314
rect 13003 28262 13055 28314
rect 13067 28262 13119 28314
rect 3792 28203 3844 28212
rect 3792 28169 3801 28203
rect 3801 28169 3835 28203
rect 3835 28169 3844 28203
rect 3792 28160 3844 28169
rect 7564 28160 7616 28212
rect 7840 28203 7892 28212
rect 7840 28169 7849 28203
rect 7849 28169 7883 28203
rect 7883 28169 7892 28203
rect 7840 28160 7892 28169
rect 5264 28092 5316 28144
rect 4252 28067 4304 28076
rect 4252 28033 4261 28067
rect 4261 28033 4295 28067
rect 4295 28033 4304 28067
rect 4252 28024 4304 28033
rect 4436 28067 4488 28076
rect 4436 28033 4445 28067
rect 4445 28033 4479 28067
rect 4479 28033 4488 28067
rect 4436 28024 4488 28033
rect 4804 28024 4856 28076
rect 4620 27956 4672 28008
rect 6092 27956 6144 28008
rect 8300 28024 8352 28076
rect 11888 28024 11940 28076
rect 12532 28160 12584 28212
rect 12716 28203 12768 28212
rect 12716 28169 12725 28203
rect 12725 28169 12759 28203
rect 12759 28169 12768 28203
rect 12716 28160 12768 28169
rect 13728 28160 13780 28212
rect 16672 28203 16724 28212
rect 16672 28169 16681 28203
rect 16681 28169 16715 28203
rect 16715 28169 16724 28203
rect 16672 28160 16724 28169
rect 13636 28092 13688 28144
rect 12440 28067 12492 28076
rect 12440 28033 12449 28067
rect 12449 28033 12483 28067
rect 12483 28033 12492 28067
rect 14280 28067 14332 28076
rect 12440 28024 12492 28033
rect 14280 28033 14298 28067
rect 14298 28033 14332 28067
rect 14280 28024 14332 28033
rect 15476 28024 15528 28076
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 7472 27956 7524 28008
rect 8208 27956 8260 28008
rect 10416 27956 10468 28008
rect 7472 27820 7524 27872
rect 8024 27863 8076 27872
rect 8024 27829 8033 27863
rect 8033 27829 8067 27863
rect 8067 27829 8076 27863
rect 8024 27820 8076 27829
rect 3915 27718 3967 27770
rect 3979 27718 4031 27770
rect 4043 27718 4095 27770
rect 4107 27718 4159 27770
rect 4171 27718 4223 27770
rect 9846 27718 9898 27770
rect 9910 27718 9962 27770
rect 9974 27718 10026 27770
rect 10038 27718 10090 27770
rect 10102 27718 10154 27770
rect 15776 27718 15828 27770
rect 15840 27718 15892 27770
rect 15904 27718 15956 27770
rect 15968 27718 16020 27770
rect 16032 27718 16084 27770
rect 5908 27659 5960 27668
rect 5908 27625 5917 27659
rect 5917 27625 5951 27659
rect 5951 27625 5960 27659
rect 5908 27616 5960 27625
rect 8300 27659 8352 27668
rect 8300 27625 8309 27659
rect 8309 27625 8343 27659
rect 8343 27625 8352 27659
rect 8300 27616 8352 27625
rect 13360 27659 13412 27668
rect 13360 27625 13369 27659
rect 13369 27625 13403 27659
rect 13403 27625 13412 27659
rect 13360 27616 13412 27625
rect 14280 27659 14332 27668
rect 14280 27625 14289 27659
rect 14289 27625 14323 27659
rect 14323 27625 14332 27659
rect 14280 27616 14332 27625
rect 9772 27548 9824 27600
rect 10416 27548 10468 27600
rect 13544 27591 13596 27600
rect 13544 27557 13553 27591
rect 13553 27557 13587 27591
rect 13587 27557 13596 27591
rect 13544 27548 13596 27557
rect 9680 27455 9732 27464
rect 9680 27421 9689 27455
rect 9689 27421 9723 27455
rect 9723 27421 9732 27455
rect 9680 27412 9732 27421
rect 10232 27480 10284 27532
rect 10324 27412 10376 27464
rect 11336 27455 11388 27464
rect 11336 27421 11345 27455
rect 11345 27421 11379 27455
rect 11379 27421 11388 27455
rect 11336 27412 11388 27421
rect 11612 27455 11664 27464
rect 11612 27421 11646 27455
rect 11646 27421 11664 27455
rect 11612 27412 11664 27421
rect 12348 27412 12400 27464
rect 14004 27412 14056 27464
rect 4436 27344 4488 27396
rect 5724 27387 5776 27396
rect 5724 27353 5733 27387
rect 5733 27353 5767 27387
rect 5767 27353 5776 27387
rect 5724 27344 5776 27353
rect 4712 27276 4764 27328
rect 5448 27276 5500 27328
rect 7288 27344 7340 27396
rect 11888 27344 11940 27396
rect 7380 27276 7432 27328
rect 9404 27319 9456 27328
rect 9404 27285 9413 27319
rect 9413 27285 9447 27319
rect 9447 27285 9456 27319
rect 9404 27276 9456 27285
rect 12256 27276 12308 27328
rect 13820 27344 13872 27396
rect 6880 27174 6932 27226
rect 6944 27174 6996 27226
rect 7008 27174 7060 27226
rect 7072 27174 7124 27226
rect 7136 27174 7188 27226
rect 12811 27174 12863 27226
rect 12875 27174 12927 27226
rect 12939 27174 12991 27226
rect 13003 27174 13055 27226
rect 13067 27174 13119 27226
rect 4712 27072 4764 27124
rect 5724 27072 5776 27124
rect 9680 27072 9732 27124
rect 11612 27072 11664 27124
rect 12440 27072 12492 27124
rect 16856 27072 16908 27124
rect 7288 27004 7340 27056
rect 9404 27047 9456 27056
rect 4528 26936 4580 26988
rect 4988 26979 5040 26988
rect 4988 26945 4997 26979
rect 4997 26945 5031 26979
rect 5031 26945 5040 26979
rect 4988 26936 5040 26945
rect 8392 26979 8444 26988
rect 9404 27013 9438 27047
rect 9438 27013 9456 27047
rect 9404 27004 9456 27013
rect 12532 27004 12584 27056
rect 13360 27004 13412 27056
rect 8392 26945 8410 26979
rect 8410 26945 8444 26979
rect 8392 26936 8444 26945
rect 9772 26936 9824 26988
rect 12072 26936 12124 26988
rect 12256 26936 12308 26988
rect 16764 26979 16816 26988
rect 16764 26945 16773 26979
rect 16773 26945 16807 26979
rect 16807 26945 16816 26979
rect 16764 26936 16816 26945
rect 16948 26936 17000 26988
rect 12624 26868 12676 26920
rect 1492 26775 1544 26784
rect 1492 26741 1501 26775
rect 1501 26741 1535 26775
rect 1535 26741 1544 26775
rect 1492 26732 1544 26741
rect 4436 26732 4488 26784
rect 7472 26800 7524 26852
rect 11704 26800 11756 26852
rect 13452 26800 13504 26852
rect 12440 26775 12492 26784
rect 12440 26741 12449 26775
rect 12449 26741 12483 26775
rect 12483 26741 12492 26775
rect 12440 26732 12492 26741
rect 3915 26630 3967 26682
rect 3979 26630 4031 26682
rect 4043 26630 4095 26682
rect 4107 26630 4159 26682
rect 4171 26630 4223 26682
rect 9846 26630 9898 26682
rect 9910 26630 9962 26682
rect 9974 26630 10026 26682
rect 10038 26630 10090 26682
rect 10102 26630 10154 26682
rect 15776 26630 15828 26682
rect 15840 26630 15892 26682
rect 15904 26630 15956 26682
rect 15968 26630 16020 26682
rect 16032 26630 16084 26682
rect 5540 26528 5592 26580
rect 1676 26460 1728 26512
rect 8024 26528 8076 26580
rect 8392 26571 8444 26580
rect 8392 26537 8401 26571
rect 8401 26537 8435 26571
rect 8435 26537 8444 26571
rect 8392 26528 8444 26537
rect 12072 26571 12124 26580
rect 12072 26537 12081 26571
rect 12081 26537 12115 26571
rect 12115 26537 12124 26571
rect 12072 26528 12124 26537
rect 3608 26392 3660 26444
rect 4436 26324 4488 26376
rect 4712 26367 4764 26376
rect 4712 26333 4721 26367
rect 4721 26333 4755 26367
rect 4755 26333 4764 26367
rect 4712 26324 4764 26333
rect 5080 26367 5132 26376
rect 5080 26333 5089 26367
rect 5089 26333 5123 26367
rect 5123 26333 5132 26367
rect 5080 26324 5132 26333
rect 7288 26392 7340 26444
rect 7380 26367 7432 26376
rect 7380 26333 7389 26367
rect 7389 26333 7423 26367
rect 7423 26333 7432 26367
rect 7380 26324 7432 26333
rect 7564 26367 7616 26376
rect 7564 26333 7573 26367
rect 7573 26333 7607 26367
rect 7607 26333 7616 26367
rect 7564 26324 7616 26333
rect 8024 26324 8076 26376
rect 8392 26367 8444 26376
rect 8392 26333 8401 26367
rect 8401 26333 8435 26367
rect 8435 26333 8444 26367
rect 8392 26324 8444 26333
rect 9772 26392 9824 26444
rect 12440 26435 12492 26444
rect 12440 26401 12449 26435
rect 12449 26401 12483 26435
rect 12483 26401 12492 26435
rect 12440 26392 12492 26401
rect 5172 26256 5224 26308
rect 6368 26256 6420 26308
rect 11704 26324 11756 26376
rect 14096 26324 14148 26376
rect 5356 26188 5408 26240
rect 10416 26256 10468 26308
rect 10692 26188 10744 26240
rect 6880 26086 6932 26138
rect 6944 26086 6996 26138
rect 7008 26086 7060 26138
rect 7072 26086 7124 26138
rect 7136 26086 7188 26138
rect 12811 26086 12863 26138
rect 12875 26086 12927 26138
rect 12939 26086 12991 26138
rect 13003 26086 13055 26138
rect 13067 26086 13119 26138
rect 6368 26027 6420 26036
rect 6368 25993 6377 26027
rect 6377 25993 6411 26027
rect 6411 25993 6420 26027
rect 6368 25984 6420 25993
rect 8392 25984 8444 26036
rect 10324 25984 10376 26036
rect 10416 25984 10468 26036
rect 12624 25984 12676 26036
rect 5632 25916 5684 25968
rect 7288 25916 7340 25968
rect 11336 25916 11388 25968
rect 3608 25891 3660 25900
rect 3608 25857 3617 25891
rect 3617 25857 3651 25891
rect 3651 25857 3660 25891
rect 3608 25848 3660 25857
rect 3700 25848 3752 25900
rect 7380 25848 7432 25900
rect 10416 25848 10468 25900
rect 10692 25891 10744 25900
rect 10692 25857 10701 25891
rect 10701 25857 10735 25891
rect 10735 25857 10744 25891
rect 10692 25848 10744 25857
rect 12808 25848 12860 25900
rect 15476 25891 15528 25900
rect 15476 25857 15485 25891
rect 15485 25857 15519 25891
rect 15519 25857 15528 25891
rect 15476 25848 15528 25857
rect 16580 25848 16632 25900
rect 6920 25780 6972 25832
rect 7564 25780 7616 25832
rect 11612 25780 11664 25832
rect 16764 25823 16816 25832
rect 16764 25789 16773 25823
rect 16773 25789 16807 25823
rect 16807 25789 16816 25823
rect 16764 25780 16816 25789
rect 5264 25712 5316 25764
rect 4988 25687 5040 25696
rect 4988 25653 4997 25687
rect 4997 25653 5031 25687
rect 5031 25653 5040 25687
rect 4988 25644 5040 25653
rect 15568 25644 15620 25696
rect 17960 25712 18012 25764
rect 17040 25687 17092 25696
rect 17040 25653 17049 25687
rect 17049 25653 17083 25687
rect 17083 25653 17092 25687
rect 17040 25644 17092 25653
rect 3915 25542 3967 25594
rect 3979 25542 4031 25594
rect 4043 25542 4095 25594
rect 4107 25542 4159 25594
rect 4171 25542 4223 25594
rect 9846 25542 9898 25594
rect 9910 25542 9962 25594
rect 9974 25542 10026 25594
rect 10038 25542 10090 25594
rect 10102 25542 10154 25594
rect 15776 25542 15828 25594
rect 15840 25542 15892 25594
rect 15904 25542 15956 25594
rect 15968 25542 16020 25594
rect 16032 25542 16084 25594
rect 3700 25440 3752 25492
rect 5264 25483 5316 25492
rect 5264 25449 5273 25483
rect 5273 25449 5307 25483
rect 5307 25449 5316 25483
rect 5264 25440 5316 25449
rect 5632 25440 5684 25492
rect 6920 25440 6972 25492
rect 12808 25440 12860 25492
rect 16672 25440 16724 25492
rect 16856 25440 16908 25492
rect 3240 25372 3292 25424
rect 3700 25236 3752 25288
rect 4988 25304 5040 25356
rect 4252 25279 4304 25288
rect 4252 25245 4261 25279
rect 4261 25245 4295 25279
rect 4295 25245 4304 25279
rect 4252 25236 4304 25245
rect 4804 25236 4856 25288
rect 5356 25236 5408 25288
rect 5724 25236 5776 25288
rect 11612 25372 11664 25424
rect 12072 25372 12124 25424
rect 16304 25372 16356 25424
rect 12256 25304 12308 25356
rect 4620 25168 4672 25220
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 12532 25279 12584 25288
rect 11796 25236 11848 25245
rect 12532 25245 12541 25279
rect 12541 25245 12575 25279
rect 12575 25245 12584 25279
rect 12532 25236 12584 25245
rect 14464 25279 14516 25288
rect 5632 25100 5684 25152
rect 11520 25168 11572 25220
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 10416 25100 10468 25152
rect 11152 25143 11204 25152
rect 11152 25109 11161 25143
rect 11161 25109 11195 25143
rect 11195 25109 11204 25143
rect 11152 25100 11204 25109
rect 11336 25100 11388 25152
rect 14832 25100 14884 25152
rect 15292 25143 15344 25152
rect 15292 25109 15301 25143
rect 15301 25109 15335 25143
rect 15335 25109 15344 25143
rect 15292 25100 15344 25109
rect 15568 25279 15620 25288
rect 15568 25245 15577 25279
rect 15577 25245 15611 25279
rect 15611 25245 15620 25279
rect 15568 25236 15620 25245
rect 16580 25304 16632 25356
rect 16672 25236 16724 25288
rect 16304 25168 16356 25220
rect 16764 25211 16816 25220
rect 16764 25177 16773 25211
rect 16773 25177 16807 25211
rect 16807 25177 16816 25211
rect 16764 25168 16816 25177
rect 17132 25100 17184 25152
rect 6880 24998 6932 25050
rect 6944 24998 6996 25050
rect 7008 24998 7060 25050
rect 7072 24998 7124 25050
rect 7136 24998 7188 25050
rect 12811 24998 12863 25050
rect 12875 24998 12927 25050
rect 12939 24998 12991 25050
rect 13003 24998 13055 25050
rect 13067 24998 13119 25050
rect 12532 24896 12584 24948
rect 14464 24896 14516 24948
rect 11152 24828 11204 24880
rect 5080 24803 5132 24812
rect 5080 24769 5089 24803
rect 5089 24769 5123 24803
rect 5123 24769 5132 24803
rect 5080 24760 5132 24769
rect 5172 24760 5224 24812
rect 5356 24760 5408 24812
rect 5632 24803 5684 24812
rect 5632 24769 5641 24803
rect 5641 24769 5675 24803
rect 5675 24769 5684 24803
rect 5632 24760 5684 24769
rect 5816 24803 5868 24812
rect 5816 24769 5825 24803
rect 5825 24769 5859 24803
rect 5859 24769 5868 24803
rect 5816 24760 5868 24769
rect 16948 24896 17000 24948
rect 15292 24760 15344 24812
rect 16672 24803 16724 24812
rect 5540 24735 5592 24744
rect 5540 24701 5549 24735
rect 5549 24701 5583 24735
rect 5583 24701 5592 24735
rect 5540 24692 5592 24701
rect 14648 24692 14700 24744
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17040 24760 17092 24812
rect 18052 24760 18104 24812
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 12256 24556 12308 24608
rect 17408 24692 17460 24744
rect 15108 24556 15160 24608
rect 17592 24556 17644 24608
rect 3915 24454 3967 24506
rect 3979 24454 4031 24506
rect 4043 24454 4095 24506
rect 4107 24454 4159 24506
rect 4171 24454 4223 24506
rect 9846 24454 9898 24506
rect 9910 24454 9962 24506
rect 9974 24454 10026 24506
rect 10038 24454 10090 24506
rect 10102 24454 10154 24506
rect 15776 24454 15828 24506
rect 15840 24454 15892 24506
rect 15904 24454 15956 24506
rect 15968 24454 16020 24506
rect 16032 24454 16084 24506
rect 5172 24395 5224 24404
rect 5172 24361 5181 24395
rect 5181 24361 5215 24395
rect 5215 24361 5224 24395
rect 5172 24352 5224 24361
rect 15476 24352 15528 24404
rect 16764 24352 16816 24404
rect 17132 24395 17184 24404
rect 17132 24361 17141 24395
rect 17141 24361 17175 24395
rect 17175 24361 17184 24395
rect 17132 24352 17184 24361
rect 2412 24216 2464 24268
rect 3884 24216 3936 24268
rect 4344 24216 4396 24268
rect 3700 24080 3752 24132
rect 14096 24148 14148 24200
rect 14464 24148 14516 24200
rect 15200 24191 15252 24200
rect 15200 24157 15209 24191
rect 15209 24157 15243 24191
rect 15243 24157 15252 24191
rect 15200 24148 15252 24157
rect 17868 24216 17920 24268
rect 18144 24148 18196 24200
rect 2964 24055 3016 24064
rect 2964 24021 2973 24055
rect 2973 24021 3007 24055
rect 3007 24021 3016 24055
rect 2964 24012 3016 24021
rect 3148 24012 3200 24064
rect 10508 24012 10560 24064
rect 11980 24012 12032 24064
rect 15568 24080 15620 24132
rect 16580 24080 16632 24132
rect 17592 24080 17644 24132
rect 18052 24080 18104 24132
rect 16120 24012 16172 24064
rect 17408 24055 17460 24064
rect 17408 24021 17417 24055
rect 17417 24021 17451 24055
rect 17451 24021 17460 24055
rect 17408 24012 17460 24021
rect 6880 23910 6932 23962
rect 6944 23910 6996 23962
rect 7008 23910 7060 23962
rect 7072 23910 7124 23962
rect 7136 23910 7188 23962
rect 12811 23910 12863 23962
rect 12875 23910 12927 23962
rect 12939 23910 12991 23962
rect 13003 23910 13055 23962
rect 13067 23910 13119 23962
rect 4252 23808 4304 23860
rect 17408 23808 17460 23860
rect 3884 23783 3936 23792
rect 3884 23749 3893 23783
rect 3893 23749 3927 23783
rect 3927 23749 3936 23783
rect 3884 23740 3936 23749
rect 12256 23740 12308 23792
rect 2964 23715 3016 23724
rect 2964 23681 2973 23715
rect 2973 23681 3007 23715
rect 3007 23681 3016 23715
rect 2964 23672 3016 23681
rect 3240 23672 3292 23724
rect 3700 23672 3752 23724
rect 7196 23715 7248 23724
rect 7196 23681 7205 23715
rect 7205 23681 7239 23715
rect 7239 23681 7248 23715
rect 7196 23672 7248 23681
rect 8208 23672 8260 23724
rect 6736 23604 6788 23656
rect 7288 23604 7340 23656
rect 13636 23604 13688 23656
rect 8116 23536 8168 23588
rect 3424 23511 3476 23520
rect 3424 23477 3433 23511
rect 3433 23477 3467 23511
rect 3467 23477 3476 23511
rect 3424 23468 3476 23477
rect 7564 23468 7616 23520
rect 7840 23511 7892 23520
rect 7840 23477 7849 23511
rect 7849 23477 7883 23511
rect 7883 23477 7892 23511
rect 7840 23468 7892 23477
rect 13268 23511 13320 23520
rect 13268 23477 13277 23511
rect 13277 23477 13311 23511
rect 13311 23477 13320 23511
rect 13268 23468 13320 23477
rect 14832 23715 14884 23724
rect 15200 23740 15252 23792
rect 14832 23681 14850 23715
rect 14850 23681 14884 23715
rect 14832 23672 14884 23681
rect 16120 23715 16172 23724
rect 16120 23681 16129 23715
rect 16129 23681 16163 23715
rect 16163 23681 16172 23715
rect 16120 23672 16172 23681
rect 16764 23715 16816 23724
rect 16764 23681 16773 23715
rect 16773 23681 16807 23715
rect 16807 23681 16816 23715
rect 16764 23672 16816 23681
rect 17592 23672 17644 23724
rect 13820 23468 13872 23520
rect 16212 23468 16264 23520
rect 3915 23366 3967 23418
rect 3979 23366 4031 23418
rect 4043 23366 4095 23418
rect 4107 23366 4159 23418
rect 4171 23366 4223 23418
rect 9846 23366 9898 23418
rect 9910 23366 9962 23418
rect 9974 23366 10026 23418
rect 10038 23366 10090 23418
rect 10102 23366 10154 23418
rect 15776 23366 15828 23418
rect 15840 23366 15892 23418
rect 15904 23366 15956 23418
rect 15968 23366 16020 23418
rect 16032 23366 16084 23418
rect 3332 23264 3384 23316
rect 3424 23264 3476 23316
rect 5724 23264 5776 23316
rect 9128 23307 9180 23316
rect 2964 23196 3016 23248
rect 3240 23128 3292 23180
rect 2872 23103 2924 23112
rect 2872 23069 2881 23103
rect 2881 23069 2915 23103
rect 2915 23069 2924 23103
rect 2872 23060 2924 23069
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 2964 23060 3016 23069
rect 3148 23103 3200 23112
rect 3148 23069 3157 23103
rect 3157 23069 3191 23103
rect 3191 23069 3200 23103
rect 3148 23060 3200 23069
rect 5632 23103 5684 23112
rect 5632 23069 5641 23103
rect 5641 23069 5675 23103
rect 5675 23069 5684 23103
rect 9128 23273 9137 23307
rect 9137 23273 9171 23307
rect 9171 23273 9180 23307
rect 9128 23264 9180 23273
rect 5632 23060 5684 23069
rect 6460 23060 6512 23112
rect 7288 23060 7340 23112
rect 8300 23103 8352 23112
rect 8300 23069 8309 23103
rect 8309 23069 8343 23103
rect 8343 23069 8352 23103
rect 8300 23060 8352 23069
rect 13636 23196 13688 23248
rect 13452 23171 13504 23180
rect 13452 23137 13461 23171
rect 13461 23137 13495 23171
rect 13495 23137 13504 23171
rect 13452 23128 13504 23137
rect 14556 23196 14608 23248
rect 16580 23128 16632 23180
rect 16764 23171 16816 23180
rect 16764 23137 16773 23171
rect 16773 23137 16807 23171
rect 16807 23137 16816 23171
rect 16764 23128 16816 23137
rect 10232 23060 10284 23112
rect 13176 23103 13228 23112
rect 13176 23069 13185 23103
rect 13185 23069 13219 23103
rect 13219 23069 13228 23103
rect 13176 23060 13228 23069
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 6092 23035 6144 23044
rect 6092 23001 6101 23035
rect 6101 23001 6135 23035
rect 6135 23001 6144 23035
rect 6092 22992 6144 23001
rect 4712 22924 4764 22976
rect 5172 22967 5224 22976
rect 5172 22933 5181 22967
rect 5181 22933 5215 22967
rect 5215 22933 5224 22967
rect 5172 22924 5224 22933
rect 6000 22924 6052 22976
rect 6368 22924 6420 22976
rect 8208 22992 8260 23044
rect 9312 23035 9364 23044
rect 8392 22967 8444 22976
rect 8392 22933 8401 22967
rect 8401 22933 8435 22967
rect 8435 22933 8444 22967
rect 8392 22924 8444 22933
rect 9312 23001 9321 23035
rect 9321 23001 9355 23035
rect 9355 23001 9364 23035
rect 9312 22992 9364 23001
rect 13820 23060 13872 23112
rect 16028 23060 16080 23112
rect 14648 22992 14700 23044
rect 17132 22992 17184 23044
rect 10508 22924 10560 22976
rect 12624 22924 12676 22976
rect 13544 22924 13596 22976
rect 16948 22924 17000 22976
rect 18052 22924 18104 22976
rect 6880 22822 6932 22874
rect 6944 22822 6996 22874
rect 7008 22822 7060 22874
rect 7072 22822 7124 22874
rect 7136 22822 7188 22874
rect 12811 22822 12863 22874
rect 12875 22822 12927 22874
rect 12939 22822 12991 22874
rect 13003 22822 13055 22874
rect 13067 22822 13119 22874
rect 3240 22763 3292 22772
rect 3240 22729 3249 22763
rect 3249 22729 3283 22763
rect 3283 22729 3292 22763
rect 3240 22720 3292 22729
rect 3792 22763 3844 22772
rect 3792 22729 3801 22763
rect 3801 22729 3835 22763
rect 3835 22729 3844 22763
rect 3792 22720 3844 22729
rect 4712 22720 4764 22772
rect 5448 22720 5500 22772
rect 6368 22720 6420 22772
rect 8300 22720 8352 22772
rect 13176 22720 13228 22772
rect 2872 22584 2924 22636
rect 3332 22584 3384 22636
rect 4436 22627 4488 22636
rect 4436 22593 4445 22627
rect 4445 22593 4479 22627
rect 4479 22593 4488 22627
rect 4436 22584 4488 22593
rect 5172 22584 5224 22636
rect 7656 22584 7708 22636
rect 8392 22652 8444 22704
rect 9128 22652 9180 22704
rect 3240 22559 3292 22568
rect 3240 22525 3249 22559
rect 3249 22525 3283 22559
rect 3283 22525 3292 22559
rect 3240 22516 3292 22525
rect 7380 22516 7432 22568
rect 8300 22516 8352 22568
rect 2964 22448 3016 22500
rect 5724 22380 5776 22432
rect 9036 22380 9088 22432
rect 9312 22380 9364 22432
rect 10508 22627 10560 22636
rect 10508 22593 10517 22627
rect 10517 22593 10551 22627
rect 10551 22593 10560 22627
rect 10508 22584 10560 22593
rect 11520 22627 11572 22636
rect 11520 22593 11529 22627
rect 11529 22593 11563 22627
rect 11563 22593 11572 22627
rect 11520 22584 11572 22593
rect 12532 22627 12584 22636
rect 12532 22593 12566 22627
rect 12566 22593 12584 22627
rect 15016 22627 15068 22636
rect 12532 22584 12584 22593
rect 15016 22593 15025 22627
rect 15025 22593 15059 22627
rect 15059 22593 15068 22627
rect 15016 22584 15068 22593
rect 15660 22584 15712 22636
rect 16028 22584 16080 22636
rect 16764 22584 16816 22636
rect 16948 22627 17000 22636
rect 16948 22593 16982 22627
rect 16982 22593 17000 22627
rect 16948 22584 17000 22593
rect 11244 22516 11296 22568
rect 12256 22559 12308 22568
rect 12256 22525 12265 22559
rect 12265 22525 12299 22559
rect 12299 22525 12308 22559
rect 12256 22516 12308 22525
rect 14556 22559 14608 22568
rect 14556 22525 14565 22559
rect 14565 22525 14599 22559
rect 14599 22525 14608 22559
rect 14556 22516 14608 22525
rect 13636 22491 13688 22500
rect 13636 22457 13645 22491
rect 13645 22457 13679 22491
rect 13679 22457 13688 22491
rect 13636 22448 13688 22457
rect 14648 22448 14700 22500
rect 11612 22380 11664 22432
rect 18144 22380 18196 22432
rect 3915 22278 3967 22330
rect 3979 22278 4031 22330
rect 4043 22278 4095 22330
rect 4107 22278 4159 22330
rect 4171 22278 4223 22330
rect 9846 22278 9898 22330
rect 9910 22278 9962 22330
rect 9974 22278 10026 22330
rect 10038 22278 10090 22330
rect 10102 22278 10154 22330
rect 15776 22278 15828 22330
rect 15840 22278 15892 22330
rect 15904 22278 15956 22330
rect 15968 22278 16020 22330
rect 16032 22278 16084 22330
rect 2780 22176 2832 22228
rect 3240 22176 3292 22228
rect 7656 22176 7708 22228
rect 13268 22176 13320 22228
rect 13360 22108 13412 22160
rect 5724 22083 5776 22092
rect 5724 22049 5733 22083
rect 5733 22049 5767 22083
rect 5767 22049 5776 22083
rect 5724 22040 5776 22049
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 10692 22040 10744 22092
rect 2780 21972 2832 22024
rect 3700 21972 3752 22024
rect 4344 21972 4396 22024
rect 4528 21972 4580 22024
rect 8300 21972 8352 22024
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 11428 22015 11480 22024
rect 9128 21972 9180 21981
rect 11428 21981 11437 22015
rect 11437 21981 11471 22015
rect 11471 21981 11480 22015
rect 11428 21972 11480 21981
rect 13452 22040 13504 22092
rect 13544 22083 13596 22092
rect 13544 22049 13553 22083
rect 13553 22049 13587 22083
rect 13587 22049 13596 22083
rect 13544 22040 13596 22049
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 15660 22040 15712 22092
rect 13268 21972 13320 21981
rect 14556 22015 14608 22024
rect 14556 21981 14565 22015
rect 14565 21981 14599 22015
rect 14599 21981 14608 22015
rect 18144 22040 18196 22092
rect 14556 21972 14608 21981
rect 2780 21836 2832 21888
rect 2964 21836 3016 21888
rect 3700 21836 3752 21888
rect 4344 21836 4396 21888
rect 5632 21836 5684 21888
rect 6736 21836 6788 21888
rect 7840 21904 7892 21956
rect 9588 21904 9640 21956
rect 13544 21904 13596 21956
rect 18052 21904 18104 21956
rect 7380 21836 7432 21888
rect 8116 21836 8168 21888
rect 8576 21836 8628 21888
rect 10968 21879 11020 21888
rect 10968 21845 10977 21879
rect 10977 21845 11011 21879
rect 11011 21845 11020 21879
rect 10968 21836 11020 21845
rect 13452 21836 13504 21888
rect 16764 21836 16816 21888
rect 17776 21836 17828 21888
rect 6880 21734 6932 21786
rect 6944 21734 6996 21786
rect 7008 21734 7060 21786
rect 7072 21734 7124 21786
rect 7136 21734 7188 21786
rect 12811 21734 12863 21786
rect 12875 21734 12927 21786
rect 12939 21734 12991 21786
rect 13003 21734 13055 21786
rect 13067 21734 13119 21786
rect 2964 21496 3016 21548
rect 3332 21496 3384 21548
rect 4620 21632 4672 21684
rect 5816 21675 5868 21684
rect 5816 21641 5825 21675
rect 5825 21641 5859 21675
rect 5859 21641 5868 21675
rect 5816 21632 5868 21641
rect 10692 21632 10744 21684
rect 12532 21632 12584 21684
rect 17132 21675 17184 21684
rect 17132 21641 17141 21675
rect 17141 21641 17175 21675
rect 17175 21641 17184 21675
rect 17132 21632 17184 21641
rect 17592 21675 17644 21684
rect 17592 21641 17601 21675
rect 17601 21641 17635 21675
rect 17635 21641 17644 21675
rect 17592 21632 17644 21641
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 4252 21539 4304 21548
rect 4252 21505 4261 21539
rect 4261 21505 4295 21539
rect 4295 21505 4304 21539
rect 4804 21564 4856 21616
rect 4252 21496 4304 21505
rect 5540 21539 5592 21548
rect 2780 21428 2832 21437
rect 4528 21428 4580 21480
rect 3700 21360 3752 21412
rect 3792 21335 3844 21344
rect 3792 21301 3801 21335
rect 3801 21301 3835 21335
rect 3835 21301 3844 21335
rect 3792 21292 3844 21301
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 5724 21496 5776 21548
rect 5816 21496 5868 21548
rect 7472 21539 7524 21548
rect 7472 21505 7490 21539
rect 7490 21505 7524 21539
rect 7472 21496 7524 21505
rect 8300 21496 8352 21548
rect 8484 21539 8536 21548
rect 8484 21505 8518 21539
rect 8518 21505 8536 21539
rect 10232 21539 10284 21548
rect 8484 21496 8536 21505
rect 10232 21505 10241 21539
rect 10241 21505 10275 21539
rect 10275 21505 10284 21539
rect 10232 21496 10284 21505
rect 11888 21496 11940 21548
rect 13452 21539 13504 21548
rect 13452 21505 13461 21539
rect 13461 21505 13495 21539
rect 13495 21505 13504 21539
rect 13452 21496 13504 21505
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 17776 21539 17828 21548
rect 17776 21505 17785 21539
rect 17785 21505 17819 21539
rect 17819 21505 17828 21539
rect 17776 21496 17828 21505
rect 9680 21428 9732 21480
rect 10968 21428 11020 21480
rect 6184 21360 6236 21412
rect 5632 21292 5684 21344
rect 9588 21335 9640 21344
rect 9588 21301 9597 21335
rect 9597 21301 9631 21335
rect 9631 21301 9640 21335
rect 9588 21292 9640 21301
rect 11336 21292 11388 21344
rect 11704 21335 11756 21344
rect 11704 21301 11713 21335
rect 11713 21301 11747 21335
rect 11747 21301 11756 21335
rect 11704 21292 11756 21301
rect 3915 21190 3967 21242
rect 3979 21190 4031 21242
rect 4043 21190 4095 21242
rect 4107 21190 4159 21242
rect 4171 21190 4223 21242
rect 9846 21190 9898 21242
rect 9910 21190 9962 21242
rect 9974 21190 10026 21242
rect 10038 21190 10090 21242
rect 10102 21190 10154 21242
rect 15776 21190 15828 21242
rect 15840 21190 15892 21242
rect 15904 21190 15956 21242
rect 15968 21190 16020 21242
rect 16032 21190 16084 21242
rect 4528 21088 4580 21140
rect 16120 21088 16172 21140
rect 6184 20995 6236 21004
rect 6184 20961 6193 20995
rect 6193 20961 6227 20995
rect 6227 20961 6236 20995
rect 6184 20952 6236 20961
rect 6460 20995 6512 21004
rect 6460 20961 6469 20995
rect 6469 20961 6503 20995
rect 6503 20961 6512 20995
rect 6460 20952 6512 20961
rect 11244 20952 11296 21004
rect 4436 20884 4488 20936
rect 7380 20884 7432 20936
rect 8116 20927 8168 20936
rect 8116 20893 8125 20927
rect 8125 20893 8159 20927
rect 8159 20893 8168 20927
rect 8116 20884 8168 20893
rect 8300 20884 8352 20936
rect 11612 20927 11664 20936
rect 11612 20893 11646 20927
rect 11646 20893 11664 20927
rect 11612 20884 11664 20893
rect 12716 20884 12768 20936
rect 13360 20927 13412 20936
rect 13360 20893 13369 20927
rect 13369 20893 13403 20927
rect 13403 20893 13412 20927
rect 13360 20884 13412 20893
rect 3792 20816 3844 20868
rect 9588 20816 9640 20868
rect 10784 20816 10836 20868
rect 7656 20791 7708 20800
rect 7656 20757 7665 20791
rect 7665 20757 7699 20791
rect 7699 20757 7708 20791
rect 7656 20748 7708 20757
rect 9496 20791 9548 20800
rect 9496 20757 9505 20791
rect 9505 20757 9539 20791
rect 9539 20757 9548 20791
rect 9496 20748 9548 20757
rect 13176 20748 13228 20800
rect 6880 20646 6932 20698
rect 6944 20646 6996 20698
rect 7008 20646 7060 20698
rect 7072 20646 7124 20698
rect 7136 20646 7188 20698
rect 12811 20646 12863 20698
rect 12875 20646 12927 20698
rect 12939 20646 12991 20698
rect 13003 20646 13055 20698
rect 13067 20646 13119 20698
rect 4252 20544 4304 20596
rect 7472 20544 7524 20596
rect 8392 20544 8444 20596
rect 8576 20544 8628 20596
rect 10232 20544 10284 20596
rect 11428 20544 11480 20596
rect 3608 20476 3660 20528
rect 3700 20451 3752 20460
rect 3700 20417 3709 20451
rect 3709 20417 3743 20451
rect 3743 20417 3752 20451
rect 3700 20408 3752 20417
rect 7656 20476 7708 20528
rect 9496 20476 9548 20528
rect 5724 20408 5776 20460
rect 6460 20408 6512 20460
rect 7380 20408 7432 20460
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 9036 20451 9088 20460
rect 7840 20408 7892 20417
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9036 20408 9088 20417
rect 11888 20476 11940 20528
rect 15292 20476 15344 20528
rect 8484 20272 8536 20324
rect 6000 20204 6052 20256
rect 8576 20204 8628 20256
rect 9680 20204 9732 20256
rect 12716 20408 12768 20460
rect 11336 20340 11388 20392
rect 12164 20315 12216 20324
rect 12164 20281 12173 20315
rect 12173 20281 12207 20315
rect 12207 20281 12216 20315
rect 12164 20272 12216 20281
rect 10232 20247 10284 20256
rect 10232 20213 10241 20247
rect 10241 20213 10275 20247
rect 10275 20213 10284 20247
rect 10232 20204 10284 20213
rect 10968 20204 11020 20256
rect 3915 20102 3967 20154
rect 3979 20102 4031 20154
rect 4043 20102 4095 20154
rect 4107 20102 4159 20154
rect 4171 20102 4223 20154
rect 9846 20102 9898 20154
rect 9910 20102 9962 20154
rect 9974 20102 10026 20154
rect 10038 20102 10090 20154
rect 10102 20102 10154 20154
rect 15776 20102 15828 20154
rect 15840 20102 15892 20154
rect 15904 20102 15956 20154
rect 15968 20102 16020 20154
rect 16032 20102 16084 20154
rect 7840 20000 7892 20052
rect 10784 20043 10836 20052
rect 10784 20009 10793 20043
rect 10793 20009 10827 20043
rect 10827 20009 10836 20043
rect 10784 20000 10836 20009
rect 10692 19932 10744 19984
rect 15016 19932 15068 19984
rect 11336 19864 11388 19916
rect 8116 19796 8168 19848
rect 9496 19796 9548 19848
rect 10968 19839 11020 19848
rect 10968 19805 10977 19839
rect 10977 19805 11011 19839
rect 11011 19805 11020 19839
rect 10968 19796 11020 19805
rect 15108 19796 15160 19848
rect 15660 19796 15712 19848
rect 12716 19728 12768 19780
rect 9496 19703 9548 19712
rect 9496 19669 9505 19703
rect 9505 19669 9539 19703
rect 9539 19669 9548 19703
rect 9496 19660 9548 19669
rect 16672 19660 16724 19712
rect 6880 19558 6932 19610
rect 6944 19558 6996 19610
rect 7008 19558 7060 19610
rect 7072 19558 7124 19610
rect 7136 19558 7188 19610
rect 12811 19558 12863 19610
rect 12875 19558 12927 19610
rect 12939 19558 12991 19610
rect 13003 19558 13055 19610
rect 13067 19558 13119 19610
rect 15200 19456 15252 19508
rect 9772 19388 9824 19440
rect 15108 19388 15160 19440
rect 9680 19320 9732 19372
rect 12716 19320 12768 19372
rect 13360 19252 13412 19304
rect 14372 19252 14424 19304
rect 13176 19116 13228 19168
rect 15016 19320 15068 19372
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 16212 19252 16264 19304
rect 15384 19184 15436 19236
rect 16120 19116 16172 19168
rect 16856 19159 16908 19168
rect 16856 19125 16865 19159
rect 16865 19125 16899 19159
rect 16899 19125 16908 19159
rect 16856 19116 16908 19125
rect 3915 19014 3967 19066
rect 3979 19014 4031 19066
rect 4043 19014 4095 19066
rect 4107 19014 4159 19066
rect 4171 19014 4223 19066
rect 9846 19014 9898 19066
rect 9910 19014 9962 19066
rect 9974 19014 10026 19066
rect 10038 19014 10090 19066
rect 10102 19014 10154 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 15904 19014 15956 19066
rect 15968 19014 16020 19066
rect 16032 19014 16084 19066
rect 5632 18955 5684 18964
rect 5632 18921 5641 18955
rect 5641 18921 5675 18955
rect 5675 18921 5684 18955
rect 5632 18912 5684 18921
rect 15108 18912 15160 18964
rect 16120 18912 16172 18964
rect 12532 18844 12584 18896
rect 13176 18819 13228 18828
rect 13176 18785 13185 18819
rect 13185 18785 13219 18819
rect 13219 18785 13228 18819
rect 13176 18776 13228 18785
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 12072 18708 12124 18760
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12440 18708 12492 18717
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 14924 18708 14976 18760
rect 16764 18708 16816 18760
rect 15476 18683 15528 18692
rect 15476 18649 15494 18683
rect 15494 18649 15528 18683
rect 15476 18640 15528 18649
rect 16856 18640 16908 18692
rect 13360 18572 13412 18624
rect 6880 18470 6932 18522
rect 6944 18470 6996 18522
rect 7008 18470 7060 18522
rect 7072 18470 7124 18522
rect 7136 18470 7188 18522
rect 12811 18470 12863 18522
rect 12875 18470 12927 18522
rect 12939 18470 12991 18522
rect 13003 18470 13055 18522
rect 13067 18470 13119 18522
rect 5540 18368 5592 18420
rect 4252 18232 4304 18284
rect 5264 18232 5316 18284
rect 8208 18368 8260 18420
rect 6368 18300 6420 18352
rect 14096 18300 14148 18352
rect 1400 18071 1452 18080
rect 1400 18037 1409 18071
rect 1409 18037 1443 18071
rect 1443 18037 1452 18071
rect 1400 18028 1452 18037
rect 5540 18071 5592 18080
rect 5540 18037 5549 18071
rect 5549 18037 5583 18071
rect 5583 18037 5592 18071
rect 5540 18028 5592 18037
rect 5816 18028 5868 18080
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 14648 18275 14700 18284
rect 14648 18241 14666 18275
rect 14666 18241 14700 18275
rect 14648 18232 14700 18241
rect 15200 18300 15252 18352
rect 14924 18275 14976 18284
rect 14924 18241 14933 18275
rect 14933 18241 14967 18275
rect 14967 18241 14976 18275
rect 14924 18232 14976 18241
rect 15292 18232 15344 18284
rect 7656 18164 7708 18216
rect 12072 18164 12124 18216
rect 7196 18096 7248 18148
rect 6920 18028 6972 18080
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 12256 18028 12308 18037
rect 14556 18028 14608 18080
rect 16212 18232 16264 18284
rect 16304 18164 16356 18216
rect 17408 18096 17460 18148
rect 15200 18028 15252 18080
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 3915 17926 3967 17978
rect 3979 17926 4031 17978
rect 4043 17926 4095 17978
rect 4107 17926 4159 17978
rect 4171 17926 4223 17978
rect 9846 17926 9898 17978
rect 9910 17926 9962 17978
rect 9974 17926 10026 17978
rect 10038 17926 10090 17978
rect 10102 17926 10154 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 15904 17926 15956 17978
rect 15968 17926 16020 17978
rect 16032 17926 16084 17978
rect 4896 17824 4948 17876
rect 7196 17867 7248 17876
rect 7196 17833 7205 17867
rect 7205 17833 7239 17867
rect 7239 17833 7248 17867
rect 7196 17824 7248 17833
rect 4620 17756 4672 17808
rect 5908 17756 5960 17808
rect 9680 17756 9732 17808
rect 10508 17756 10560 17808
rect 6184 17731 6236 17740
rect 6184 17697 6193 17731
rect 6193 17697 6227 17731
rect 6227 17697 6236 17731
rect 6184 17688 6236 17697
rect 6736 17688 6788 17740
rect 7564 17688 7616 17740
rect 11520 17824 11572 17876
rect 12624 17824 12676 17876
rect 15108 17824 15160 17876
rect 11796 17756 11848 17808
rect 12716 17756 12768 17808
rect 15384 17756 15436 17808
rect 4712 17620 4764 17672
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 6276 17663 6328 17672
rect 6276 17629 6285 17663
rect 6285 17629 6319 17663
rect 6319 17629 6328 17663
rect 6276 17620 6328 17629
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 9680 17620 9732 17672
rect 10968 17620 11020 17672
rect 7380 17595 7432 17604
rect 7380 17561 7389 17595
rect 7389 17561 7423 17595
rect 7423 17561 7432 17595
rect 7380 17552 7432 17561
rect 7748 17552 7800 17604
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 6644 17484 6696 17493
rect 9864 17527 9916 17536
rect 9864 17493 9873 17527
rect 9873 17493 9907 17527
rect 9907 17493 9916 17527
rect 9864 17484 9916 17493
rect 11152 17552 11204 17604
rect 12256 17688 12308 17740
rect 11704 17663 11756 17672
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 12532 17620 12584 17672
rect 12348 17552 12400 17604
rect 12808 17663 12860 17672
rect 12808 17629 12817 17663
rect 12817 17629 12851 17663
rect 12851 17629 12860 17663
rect 13360 17663 13412 17672
rect 12808 17620 12860 17629
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 14832 17552 14884 17604
rect 16212 17688 16264 17740
rect 16396 17688 16448 17740
rect 16120 17620 16172 17672
rect 16304 17595 16356 17604
rect 16304 17561 16313 17595
rect 16313 17561 16347 17595
rect 16347 17561 16356 17595
rect 16304 17552 16356 17561
rect 15936 17527 15988 17536
rect 15936 17493 15945 17527
rect 15945 17493 15979 17527
rect 15979 17493 15988 17527
rect 15936 17484 15988 17493
rect 16120 17527 16172 17536
rect 16120 17493 16147 17527
rect 16147 17493 16172 17527
rect 16120 17484 16172 17493
rect 17592 17527 17644 17536
rect 17592 17493 17601 17527
rect 17601 17493 17635 17527
rect 17635 17493 17644 17527
rect 17592 17484 17644 17493
rect 6880 17382 6932 17434
rect 6944 17382 6996 17434
rect 7008 17382 7060 17434
rect 7072 17382 7124 17434
rect 7136 17382 7188 17434
rect 12811 17382 12863 17434
rect 12875 17382 12927 17434
rect 12939 17382 12991 17434
rect 13003 17382 13055 17434
rect 13067 17382 13119 17434
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 4620 17280 4672 17332
rect 5172 17280 5224 17332
rect 14648 17280 14700 17332
rect 15476 17280 15528 17332
rect 5540 17212 5592 17264
rect 6644 17255 6696 17264
rect 6644 17221 6678 17255
rect 6678 17221 6696 17255
rect 6644 17212 6696 17221
rect 12348 17212 12400 17264
rect 5172 17187 5224 17196
rect 3608 17076 3660 17128
rect 5172 17153 5181 17187
rect 5181 17153 5215 17187
rect 5215 17153 5224 17187
rect 5172 17144 5224 17153
rect 4620 17076 4672 17128
rect 8208 17187 8260 17196
rect 8208 17153 8217 17187
rect 8217 17153 8251 17187
rect 8251 17153 8260 17187
rect 8208 17144 8260 17153
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 8576 17187 8628 17196
rect 8576 17153 8585 17187
rect 8585 17153 8619 17187
rect 8619 17153 8628 17187
rect 8576 17144 8628 17153
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 10232 17144 10284 17196
rect 11796 17187 11848 17196
rect 5448 17119 5500 17128
rect 5448 17085 5457 17119
rect 5457 17085 5491 17119
rect 5491 17085 5500 17119
rect 5448 17076 5500 17085
rect 3792 17008 3844 17060
rect 7380 17076 7432 17128
rect 10692 17076 10744 17128
rect 4252 16940 4304 16992
rect 4344 16940 4396 16992
rect 11152 17008 11204 17060
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 11704 17076 11756 17128
rect 12256 17144 12308 17196
rect 13452 17144 13504 17196
rect 13268 17076 13320 17128
rect 15936 17212 15988 17264
rect 14832 17187 14884 17196
rect 14832 17153 14841 17187
rect 14841 17153 14875 17187
rect 14875 17153 14884 17187
rect 14832 17144 14884 17153
rect 15200 17144 15252 17196
rect 16672 17280 16724 17332
rect 17960 17280 18012 17332
rect 16764 17144 16816 17196
rect 17316 17144 17368 17196
rect 16028 17076 16080 17128
rect 12256 17008 12308 17060
rect 12716 17051 12768 17060
rect 12716 17017 12725 17051
rect 12725 17017 12759 17051
rect 12759 17017 12768 17051
rect 12716 17008 12768 17017
rect 13452 17008 13504 17060
rect 7012 16940 7064 16992
rect 8024 16940 8076 16992
rect 8944 16983 8996 16992
rect 8944 16949 8953 16983
rect 8953 16949 8987 16983
rect 8987 16949 8996 16983
rect 8944 16940 8996 16949
rect 9680 16983 9732 16992
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 12624 16940 12676 16992
rect 15016 16940 15068 16992
rect 3915 16838 3967 16890
rect 3979 16838 4031 16890
rect 4043 16838 4095 16890
rect 4107 16838 4159 16890
rect 4171 16838 4223 16890
rect 9846 16838 9898 16890
rect 9910 16838 9962 16890
rect 9974 16838 10026 16890
rect 10038 16838 10090 16890
rect 10102 16838 10154 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 15904 16838 15956 16890
rect 15968 16838 16020 16890
rect 16032 16838 16084 16890
rect 5172 16736 5224 16788
rect 7012 16736 7064 16788
rect 8300 16736 8352 16788
rect 10692 16779 10744 16788
rect 6276 16668 6328 16720
rect 3516 16532 3568 16584
rect 3332 16464 3384 16516
rect 3792 16532 3844 16584
rect 4344 16575 4396 16584
rect 4344 16541 4378 16575
rect 4378 16541 4396 16575
rect 4344 16532 4396 16541
rect 10692 16745 10701 16779
rect 10701 16745 10735 16779
rect 10735 16745 10744 16779
rect 10692 16736 10744 16745
rect 11244 16736 11296 16788
rect 12348 16736 12400 16788
rect 14096 16736 14148 16788
rect 16764 16736 16816 16788
rect 12256 16668 12308 16720
rect 13268 16711 13320 16720
rect 13268 16677 13277 16711
rect 13277 16677 13311 16711
rect 13311 16677 13320 16711
rect 13268 16668 13320 16677
rect 7012 16643 7064 16652
rect 7012 16609 7021 16643
rect 7021 16609 7055 16643
rect 7055 16609 7064 16643
rect 7012 16600 7064 16609
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 13452 16600 13504 16652
rect 4896 16464 4948 16516
rect 4160 16396 4212 16448
rect 5724 16396 5776 16448
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 7564 16532 7616 16584
rect 8760 16532 8812 16584
rect 10140 16532 10192 16584
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 17592 16532 17644 16584
rect 9680 16464 9732 16516
rect 11888 16464 11940 16516
rect 14372 16464 14424 16516
rect 7380 16396 7432 16448
rect 12440 16396 12492 16448
rect 14832 16439 14884 16448
rect 14832 16405 14841 16439
rect 14841 16405 14875 16439
rect 14875 16405 14884 16439
rect 14832 16396 14884 16405
rect 16304 16396 16356 16448
rect 6880 16294 6932 16346
rect 6944 16294 6996 16346
rect 7008 16294 7060 16346
rect 7072 16294 7124 16346
rect 7136 16294 7188 16346
rect 12811 16294 12863 16346
rect 12875 16294 12927 16346
rect 12939 16294 12991 16346
rect 13003 16294 13055 16346
rect 13067 16294 13119 16346
rect 2964 16192 3016 16244
rect 6736 16235 6788 16244
rect 6736 16201 6745 16235
rect 6745 16201 6779 16235
rect 6779 16201 6788 16235
rect 6736 16192 6788 16201
rect 8576 16192 8628 16244
rect 10968 16235 11020 16244
rect 2780 16167 2832 16176
rect 2780 16133 2805 16167
rect 2805 16133 2832 16167
rect 2780 16124 2832 16133
rect 6184 16124 6236 16176
rect 3240 16056 3292 16108
rect 4160 16056 4212 16108
rect 5448 16056 5500 16108
rect 5724 16056 5776 16108
rect 7288 16124 7340 16176
rect 7840 16124 7892 16176
rect 8116 16124 8168 16176
rect 8024 16099 8076 16108
rect 8024 16065 8033 16099
rect 8033 16065 8067 16099
rect 8067 16065 8076 16099
rect 9680 16124 9732 16176
rect 10968 16201 10977 16235
rect 10977 16201 11011 16235
rect 11011 16201 11020 16235
rect 10968 16192 11020 16201
rect 12072 16192 12124 16244
rect 17316 16235 17368 16244
rect 17316 16201 17325 16235
rect 17325 16201 17359 16235
rect 17359 16201 17368 16235
rect 17316 16192 17368 16201
rect 10232 16124 10284 16176
rect 8024 16056 8076 16065
rect 9772 16099 9824 16108
rect 3056 15988 3108 16040
rect 3700 15988 3752 16040
rect 9772 16065 9781 16099
rect 9781 16065 9815 16099
rect 9815 16065 9824 16099
rect 9772 16056 9824 16065
rect 10140 16099 10192 16108
rect 10140 16065 10149 16099
rect 10149 16065 10183 16099
rect 10183 16065 10192 16099
rect 10140 16056 10192 16065
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 12348 16124 12400 16176
rect 10416 15988 10468 16040
rect 17500 16099 17552 16108
rect 17500 16065 17509 16099
rect 17509 16065 17543 16099
rect 17543 16065 17552 16099
rect 17500 16056 17552 16065
rect 14832 15988 14884 16040
rect 3332 15920 3384 15972
rect 6092 15920 6144 15972
rect 3424 15852 3476 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 8392 15852 8444 15904
rect 9588 15895 9640 15904
rect 9588 15861 9597 15895
rect 9597 15861 9631 15895
rect 9631 15861 9640 15895
rect 9588 15852 9640 15861
rect 3915 15750 3967 15802
rect 3979 15750 4031 15802
rect 4043 15750 4095 15802
rect 4107 15750 4159 15802
rect 4171 15750 4223 15802
rect 9846 15750 9898 15802
rect 9910 15750 9962 15802
rect 9974 15750 10026 15802
rect 10038 15750 10090 15802
rect 10102 15750 10154 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 15904 15750 15956 15802
rect 15968 15750 16020 15802
rect 16032 15750 16084 15802
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 6460 15648 6512 15700
rect 8208 15648 8260 15700
rect 10968 15648 11020 15700
rect 3332 15580 3384 15632
rect 3792 15512 3844 15564
rect 2780 15444 2832 15496
rect 3700 15444 3752 15496
rect 7656 15580 7708 15632
rect 6552 15555 6604 15564
rect 6552 15521 6561 15555
rect 6561 15521 6595 15555
rect 6595 15521 6604 15555
rect 6552 15512 6604 15521
rect 7288 15512 7340 15564
rect 6184 15444 6236 15496
rect 8300 15580 8352 15632
rect 8024 15512 8076 15564
rect 11244 15512 11296 15564
rect 11336 15512 11388 15564
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 8392 15444 8444 15453
rect 3240 15419 3292 15428
rect 3240 15385 3249 15419
rect 3249 15385 3283 15419
rect 3283 15385 3292 15419
rect 3240 15376 3292 15385
rect 4252 15376 4304 15428
rect 6092 15419 6144 15428
rect 6092 15385 6101 15419
rect 6101 15385 6135 15419
rect 6135 15385 6144 15419
rect 6092 15376 6144 15385
rect 7380 15376 7432 15428
rect 8116 15419 8168 15428
rect 8116 15385 8125 15419
rect 8125 15385 8159 15419
rect 8159 15385 8168 15419
rect 8116 15376 8168 15385
rect 10876 15376 10928 15428
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 6736 15308 6788 15360
rect 10324 15308 10376 15360
rect 12532 15444 12584 15496
rect 12072 15376 12124 15428
rect 14372 15419 14424 15428
rect 14372 15385 14381 15419
rect 14381 15385 14415 15419
rect 14415 15385 14424 15419
rect 14372 15376 14424 15385
rect 11704 15351 11756 15360
rect 11704 15317 11713 15351
rect 11713 15317 11747 15351
rect 11747 15317 11756 15351
rect 11704 15308 11756 15317
rect 11888 15308 11940 15360
rect 6880 15206 6932 15258
rect 6944 15206 6996 15258
rect 7008 15206 7060 15258
rect 7072 15206 7124 15258
rect 7136 15206 7188 15258
rect 12811 15206 12863 15258
rect 12875 15206 12927 15258
rect 12939 15206 12991 15258
rect 13003 15206 13055 15258
rect 13067 15206 13119 15258
rect 3608 15147 3660 15156
rect 3608 15113 3617 15147
rect 3617 15113 3651 15147
rect 3651 15113 3660 15147
rect 3608 15104 3660 15113
rect 3700 15104 3752 15156
rect 6552 15104 6604 15156
rect 10232 15104 10284 15156
rect 10876 15147 10928 15156
rect 10876 15113 10885 15147
rect 10885 15113 10919 15147
rect 10919 15113 10928 15147
rect 10876 15104 10928 15113
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 4252 15079 4304 15088
rect 4252 15045 4261 15079
rect 4261 15045 4295 15079
rect 4295 15045 4304 15079
rect 4252 15036 4304 15045
rect 5264 15036 5316 15088
rect 8392 15036 8444 15088
rect 3332 15011 3384 15020
rect 3332 14977 3341 15011
rect 3341 14977 3375 15011
rect 3375 14977 3384 15011
rect 3332 14968 3384 14977
rect 3424 15011 3476 15020
rect 3424 14977 3433 15011
rect 3433 14977 3467 15011
rect 3467 14977 3476 15011
rect 4436 15011 4488 15020
rect 3424 14968 3476 14977
rect 4436 14977 4445 15011
rect 4445 14977 4479 15011
rect 4479 14977 4488 15011
rect 4436 14968 4488 14977
rect 6920 15011 6972 15020
rect 6920 14977 6929 15011
rect 6929 14977 6963 15011
rect 6963 14977 6972 15011
rect 6920 14968 6972 14977
rect 7380 14968 7432 15020
rect 7748 15011 7800 15020
rect 7748 14977 7757 15011
rect 7757 14977 7791 15011
rect 7791 14977 7800 15011
rect 7748 14968 7800 14977
rect 8576 15011 8628 15020
rect 8576 14977 8585 15011
rect 8585 14977 8619 15011
rect 8619 14977 8628 15011
rect 8576 14968 8628 14977
rect 9680 15036 9732 15088
rect 10324 15079 10376 15088
rect 10324 15045 10333 15079
rect 10333 15045 10367 15079
rect 10367 15045 10376 15079
rect 10324 15036 10376 15045
rect 11980 15079 12032 15088
rect 11980 15045 11989 15079
rect 11989 15045 12023 15079
rect 12023 15045 12032 15079
rect 11980 15036 12032 15045
rect 9772 14968 9824 15020
rect 10232 14968 10284 15020
rect 11704 14968 11756 15020
rect 17960 14968 18012 15020
rect 3516 14900 3568 14952
rect 9220 14900 9272 14952
rect 9496 14900 9548 14952
rect 17868 14943 17920 14952
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 7656 14832 7708 14884
rect 10232 14832 10284 14884
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 10692 14764 10744 14816
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 3915 14662 3967 14714
rect 3979 14662 4031 14714
rect 4043 14662 4095 14714
rect 4107 14662 4159 14714
rect 4171 14662 4223 14714
rect 9846 14662 9898 14714
rect 9910 14662 9962 14714
rect 9974 14662 10026 14714
rect 10038 14662 10090 14714
rect 10102 14662 10154 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 15904 14662 15956 14714
rect 15968 14662 16020 14714
rect 16032 14662 16084 14714
rect 3056 14560 3108 14612
rect 8944 14560 8996 14612
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 6920 14492 6972 14544
rect 7840 14492 7892 14544
rect 13544 14492 13596 14544
rect 9588 14424 9640 14476
rect 4252 14356 4304 14408
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 4436 14288 4488 14340
rect 11520 14424 11572 14476
rect 10692 14356 10744 14408
rect 15568 14356 15620 14408
rect 18144 14399 18196 14408
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 9864 14331 9916 14340
rect 9864 14297 9873 14331
rect 9873 14297 9907 14331
rect 9907 14297 9916 14331
rect 9864 14288 9916 14297
rect 12072 14288 12124 14340
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 9680 14220 9732 14272
rect 15016 14220 15068 14272
rect 6880 14118 6932 14170
rect 6944 14118 6996 14170
rect 7008 14118 7060 14170
rect 7072 14118 7124 14170
rect 7136 14118 7188 14170
rect 12811 14118 12863 14170
rect 12875 14118 12927 14170
rect 12939 14118 12991 14170
rect 13003 14118 13055 14170
rect 13067 14118 13119 14170
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 9312 13948 9364 14000
rect 9864 13948 9916 14000
rect 14372 13948 14424 14000
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 16396 13880 16448 13932
rect 13360 13812 13412 13864
rect 14464 13812 14516 13864
rect 15660 13812 15712 13864
rect 14740 13787 14792 13796
rect 14740 13753 14749 13787
rect 14749 13753 14783 13787
rect 14783 13753 14792 13787
rect 14740 13744 14792 13753
rect 3915 13574 3967 13626
rect 3979 13574 4031 13626
rect 4043 13574 4095 13626
rect 4107 13574 4159 13626
rect 4171 13574 4223 13626
rect 9846 13574 9898 13626
rect 9910 13574 9962 13626
rect 9974 13574 10026 13626
rect 10038 13574 10090 13626
rect 10102 13574 10154 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 15904 13574 15956 13626
rect 15968 13574 16020 13626
rect 16032 13574 16084 13626
rect 16120 13472 16172 13524
rect 16304 13472 16356 13524
rect 17408 13515 17460 13524
rect 17408 13481 17417 13515
rect 17417 13481 17451 13515
rect 17451 13481 17460 13515
rect 17408 13472 17460 13481
rect 16212 13336 16264 13388
rect 13544 13268 13596 13320
rect 13820 13268 13872 13320
rect 14740 13268 14792 13320
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 16672 13268 16724 13320
rect 13452 13200 13504 13252
rect 14648 13200 14700 13252
rect 15660 13200 15712 13252
rect 13820 13132 13872 13184
rect 14096 13175 14148 13184
rect 14096 13141 14105 13175
rect 14105 13141 14139 13175
rect 14139 13141 14148 13175
rect 14096 13132 14148 13141
rect 16212 13175 16264 13184
rect 16212 13141 16221 13175
rect 16221 13141 16255 13175
rect 16255 13141 16264 13175
rect 16212 13132 16264 13141
rect 6880 13030 6932 13082
rect 6944 13030 6996 13082
rect 7008 13030 7060 13082
rect 7072 13030 7124 13082
rect 7136 13030 7188 13082
rect 12811 13030 12863 13082
rect 12875 13030 12927 13082
rect 12939 13030 12991 13082
rect 13003 13030 13055 13082
rect 13067 13030 13119 13082
rect 13268 12928 13320 12980
rect 8576 12903 8628 12912
rect 8576 12869 8585 12903
rect 8585 12869 8619 12903
rect 8619 12869 8628 12903
rect 8576 12860 8628 12869
rect 9772 12860 9824 12912
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 13728 12792 13780 12844
rect 14280 12792 14332 12844
rect 14740 12792 14792 12844
rect 16396 12792 16448 12844
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 16304 12724 16356 12776
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 8668 12631 8720 12640
rect 8668 12597 8677 12631
rect 8677 12597 8711 12631
rect 8711 12597 8720 12631
rect 8668 12588 8720 12597
rect 9588 12588 9640 12640
rect 9772 12588 9824 12640
rect 13360 12588 13412 12640
rect 17408 12588 17460 12640
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 3915 12486 3967 12538
rect 3979 12486 4031 12538
rect 4043 12486 4095 12538
rect 4107 12486 4159 12538
rect 4171 12486 4223 12538
rect 9846 12486 9898 12538
rect 9910 12486 9962 12538
rect 9974 12486 10026 12538
rect 10038 12486 10090 12538
rect 10102 12486 10154 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 15904 12486 15956 12538
rect 15968 12486 16020 12538
rect 16032 12486 16084 12538
rect 8576 12384 8628 12436
rect 12716 12384 12768 12436
rect 13728 12384 13780 12436
rect 14188 12384 14240 12436
rect 9036 12316 9088 12368
rect 9588 12248 9640 12300
rect 3792 12180 3844 12232
rect 8852 12180 8904 12232
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 7288 12155 7340 12164
rect 7288 12121 7322 12155
rect 7322 12121 7340 12155
rect 7288 12112 7340 12121
rect 8668 12112 8720 12164
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9772 12180 9824 12232
rect 10140 12180 10192 12232
rect 12164 12248 12216 12300
rect 14188 12248 14240 12300
rect 11612 12180 11664 12232
rect 14096 12180 14148 12232
rect 16672 12384 16724 12436
rect 14740 12316 14792 12368
rect 9312 12155 9364 12164
rect 9312 12121 9321 12155
rect 9321 12121 9355 12155
rect 9355 12121 9364 12155
rect 9312 12112 9364 12121
rect 10508 12112 10560 12164
rect 11796 12112 11848 12164
rect 13452 12112 13504 12164
rect 9680 12044 9732 12096
rect 10324 12044 10376 12096
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 14832 12180 14884 12232
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 14556 12155 14608 12164
rect 14556 12121 14591 12155
rect 14591 12121 14608 12155
rect 14556 12112 14608 12121
rect 17500 12112 17552 12164
rect 14832 12044 14884 12096
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 6880 11942 6932 11994
rect 6944 11942 6996 11994
rect 7008 11942 7060 11994
rect 7072 11942 7124 11994
rect 7136 11942 7188 11994
rect 12811 11942 12863 11994
rect 12875 11942 12927 11994
rect 12939 11942 12991 11994
rect 13003 11942 13055 11994
rect 13067 11942 13119 11994
rect 7288 11840 7340 11892
rect 9956 11840 10008 11892
rect 10508 11840 10560 11892
rect 14556 11840 14608 11892
rect 16212 11840 16264 11892
rect 7104 11772 7156 11824
rect 4988 11704 5040 11756
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5540 11747 5592 11756
rect 5080 11704 5132 11713
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 5908 11704 5960 11756
rect 8668 11772 8720 11824
rect 9220 11772 9272 11824
rect 9864 11815 9916 11824
rect 6276 11568 6328 11620
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 9036 11704 9088 11756
rect 9588 11747 9640 11756
rect 9588 11713 9597 11747
rect 9597 11713 9631 11747
rect 9631 11713 9640 11747
rect 9588 11704 9640 11713
rect 9864 11781 9873 11815
rect 9873 11781 9907 11815
rect 9907 11781 9916 11815
rect 9864 11772 9916 11781
rect 10232 11772 10284 11824
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 15016 11815 15068 11824
rect 15016 11781 15050 11815
rect 15050 11781 15068 11815
rect 15016 11772 15068 11781
rect 10324 11636 10376 11688
rect 11612 11704 11664 11756
rect 12716 11704 12768 11756
rect 14188 11704 14240 11756
rect 14556 11704 14608 11756
rect 14004 11636 14056 11688
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 8024 11568 8076 11620
rect 10140 11568 10192 11620
rect 4436 11500 4488 11552
rect 5632 11500 5684 11552
rect 7104 11500 7156 11552
rect 7932 11500 7984 11552
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 11520 11500 11572 11552
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 3915 11398 3967 11450
rect 3979 11398 4031 11450
rect 4043 11398 4095 11450
rect 4107 11398 4159 11450
rect 4171 11398 4223 11450
rect 9846 11398 9898 11450
rect 9910 11398 9962 11450
rect 9974 11398 10026 11450
rect 10038 11398 10090 11450
rect 10102 11398 10154 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 15904 11398 15956 11450
rect 15968 11398 16020 11450
rect 16032 11398 16084 11450
rect 7380 11296 7432 11348
rect 10324 11296 10376 11348
rect 11428 11296 11480 11348
rect 13176 11296 13228 11348
rect 13728 11296 13780 11348
rect 14556 11339 14608 11348
rect 14556 11305 14565 11339
rect 14565 11305 14599 11339
rect 14599 11305 14608 11339
rect 14556 11296 14608 11305
rect 15660 11296 15712 11348
rect 4988 11228 5040 11280
rect 6276 11203 6328 11212
rect 6276 11169 6285 11203
rect 6285 11169 6319 11203
rect 6319 11169 6328 11203
rect 6276 11160 6328 11169
rect 3792 11092 3844 11144
rect 7380 11160 7432 11212
rect 15476 11228 15528 11280
rect 7656 11203 7708 11212
rect 7656 11169 7665 11203
rect 7665 11169 7699 11203
rect 7699 11169 7708 11203
rect 7656 11160 7708 11169
rect 8852 11160 8904 11212
rect 11152 11160 11204 11212
rect 12072 11160 12124 11212
rect 4252 11067 4304 11076
rect 4252 11033 4286 11067
rect 4286 11033 4304 11067
rect 4252 11024 4304 11033
rect 5080 11024 5132 11076
rect 5816 10999 5868 11008
rect 5816 10965 5825 10999
rect 5825 10965 5859 10999
rect 5859 10965 5868 10999
rect 5816 10956 5868 10965
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8668 11092 8720 11144
rect 7288 11024 7340 11076
rect 7380 11024 7432 11076
rect 13544 11160 13596 11212
rect 14096 11160 14148 11212
rect 13452 11092 13504 11144
rect 14740 11092 14792 11144
rect 13360 11024 13412 11076
rect 17224 11024 17276 11076
rect 7748 10956 7800 11008
rect 9312 10956 9364 11008
rect 11520 10999 11572 11008
rect 11520 10965 11545 10999
rect 11545 10965 11572 10999
rect 11520 10956 11572 10965
rect 6880 10854 6932 10906
rect 6944 10854 6996 10906
rect 7008 10854 7060 10906
rect 7072 10854 7124 10906
rect 7136 10854 7188 10906
rect 12811 10854 12863 10906
rect 12875 10854 12927 10906
rect 12939 10854 12991 10906
rect 13003 10854 13055 10906
rect 13067 10854 13119 10906
rect 4252 10727 4304 10736
rect 4252 10693 4261 10727
rect 4261 10693 4295 10727
rect 4295 10693 4304 10727
rect 4252 10684 4304 10693
rect 7932 10752 7984 10804
rect 9588 10752 9640 10804
rect 10416 10752 10468 10804
rect 11428 10752 11480 10804
rect 14280 10752 14332 10804
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 7656 10727 7708 10736
rect 7656 10693 7665 10727
rect 7665 10693 7699 10727
rect 7699 10693 7708 10727
rect 7656 10684 7708 10693
rect 7748 10684 7800 10736
rect 4436 10659 4488 10668
rect 4436 10625 4445 10659
rect 4445 10625 4479 10659
rect 4479 10625 4488 10659
rect 4436 10616 4488 10625
rect 4804 10616 4856 10668
rect 5816 10616 5868 10668
rect 5908 10616 5960 10668
rect 8208 10616 8260 10668
rect 9312 10684 9364 10736
rect 5632 10591 5684 10600
rect 5632 10557 5641 10591
rect 5641 10557 5675 10591
rect 5675 10557 5684 10591
rect 5632 10548 5684 10557
rect 6276 10548 6328 10600
rect 9220 10616 9272 10668
rect 9772 10684 9824 10736
rect 12072 10684 12124 10736
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 10324 10616 10376 10668
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 13544 10616 13596 10668
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 4620 10480 4672 10532
rect 6000 10480 6052 10532
rect 7012 10480 7064 10532
rect 7288 10480 7340 10532
rect 10232 10548 10284 10600
rect 10600 10548 10652 10600
rect 12532 10548 12584 10600
rect 13728 10548 13780 10600
rect 7656 10412 7708 10464
rect 10508 10412 10560 10464
rect 12900 10412 12952 10464
rect 3915 10310 3967 10362
rect 3979 10310 4031 10362
rect 4043 10310 4095 10362
rect 4107 10310 4159 10362
rect 4171 10310 4223 10362
rect 9846 10310 9898 10362
rect 9910 10310 9962 10362
rect 9974 10310 10026 10362
rect 10038 10310 10090 10362
rect 10102 10310 10154 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 15904 10310 15956 10362
rect 15968 10310 16020 10362
rect 16032 10310 16084 10362
rect 5908 10208 5960 10260
rect 5816 10140 5868 10192
rect 7012 10208 7064 10260
rect 11796 10208 11848 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 7288 10140 7340 10192
rect 5540 10072 5592 10124
rect 6276 10072 6328 10124
rect 6644 10072 6696 10124
rect 7656 10072 7708 10124
rect 12164 10072 12216 10124
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 8392 10004 8444 10056
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 11980 10004 12032 10056
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 7748 9936 7800 9988
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 7380 9868 7432 9920
rect 6880 9766 6932 9818
rect 6944 9766 6996 9818
rect 7008 9766 7060 9818
rect 7072 9766 7124 9818
rect 7136 9766 7188 9818
rect 12811 9766 12863 9818
rect 12875 9766 12927 9818
rect 12939 9766 12991 9818
rect 13003 9766 13055 9818
rect 13067 9766 13119 9818
rect 12532 9664 12584 9716
rect 17500 9664 17552 9716
rect 17868 9664 17920 9716
rect 5540 9596 5592 9648
rect 6644 9639 6696 9648
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 6644 9596 6696 9605
rect 6736 9596 6788 9648
rect 7748 9639 7800 9648
rect 7748 9605 7757 9639
rect 7757 9605 7791 9639
rect 7791 9605 7800 9639
rect 7748 9596 7800 9605
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 5264 9460 5316 9512
rect 10508 9596 10560 9648
rect 8852 9528 8904 9580
rect 10232 9528 10284 9580
rect 7656 9392 7708 9444
rect 4712 9324 4764 9376
rect 10692 9324 10744 9376
rect 3915 9222 3967 9274
rect 3979 9222 4031 9274
rect 4043 9222 4095 9274
rect 4107 9222 4159 9274
rect 4171 9222 4223 9274
rect 9846 9222 9898 9274
rect 9910 9222 9962 9274
rect 9974 9222 10026 9274
rect 10038 9222 10090 9274
rect 10102 9222 10154 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 15904 9222 15956 9274
rect 15968 9222 16020 9274
rect 16032 9222 16084 9274
rect 4712 9163 4764 9172
rect 4712 9129 4721 9163
rect 4721 9129 4755 9163
rect 4755 9129 4764 9163
rect 4712 9120 4764 9129
rect 10232 9163 10284 9172
rect 10232 9129 10241 9163
rect 10241 9129 10275 9163
rect 10275 9129 10284 9163
rect 10232 9120 10284 9129
rect 11428 9120 11480 9172
rect 8024 9052 8076 9104
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 10508 8984 10560 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 6552 8959 6604 8968
rect 4804 8916 4856 8925
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 7840 8916 7892 8968
rect 8208 8916 8260 8968
rect 10416 8959 10468 8968
rect 10416 8925 10425 8959
rect 10425 8925 10459 8959
rect 10459 8925 10468 8959
rect 10416 8916 10468 8925
rect 10692 8916 10744 8968
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 11888 8916 11940 8968
rect 4528 8891 4580 8900
rect 4528 8857 4537 8891
rect 4537 8857 4571 8891
rect 4571 8857 4580 8891
rect 4528 8848 4580 8857
rect 4988 8891 5040 8900
rect 4988 8857 4997 8891
rect 4997 8857 5031 8891
rect 5031 8857 5040 8891
rect 4988 8848 5040 8857
rect 6880 8678 6932 8730
rect 6944 8678 6996 8730
rect 7008 8678 7060 8730
rect 7072 8678 7124 8730
rect 7136 8678 7188 8730
rect 12811 8678 12863 8730
rect 12875 8678 12927 8730
rect 12939 8678 12991 8730
rect 13003 8678 13055 8730
rect 13067 8678 13119 8730
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 11980 8576 12032 8628
rect 4528 8508 4580 8560
rect 3792 8440 3844 8492
rect 7380 8440 7432 8492
rect 7840 8440 7892 8492
rect 10968 8440 11020 8492
rect 8024 8415 8076 8424
rect 8024 8381 8033 8415
rect 8033 8381 8067 8415
rect 8067 8381 8076 8415
rect 8024 8372 8076 8381
rect 10508 8372 10560 8424
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 11980 8440 12032 8492
rect 13176 8440 13228 8492
rect 14648 8372 14700 8424
rect 7932 8347 7984 8356
rect 7932 8313 7941 8347
rect 7941 8313 7975 8347
rect 7975 8313 7984 8347
rect 7932 8304 7984 8313
rect 10692 8304 10744 8356
rect 7748 8236 7800 8288
rect 14096 8279 14148 8288
rect 14096 8245 14105 8279
rect 14105 8245 14139 8279
rect 14139 8245 14148 8279
rect 14096 8236 14148 8245
rect 3915 8134 3967 8186
rect 3979 8134 4031 8186
rect 4043 8134 4095 8186
rect 4107 8134 4159 8186
rect 4171 8134 4223 8186
rect 9846 8134 9898 8186
rect 9910 8134 9962 8186
rect 9974 8134 10026 8186
rect 10038 8134 10090 8186
rect 10102 8134 10154 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 15904 8134 15956 8186
rect 15968 8134 16020 8186
rect 16032 8134 16084 8186
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 14188 8032 14240 8084
rect 14924 8075 14976 8084
rect 14924 8041 14933 8075
rect 14933 8041 14967 8075
rect 14967 8041 14976 8075
rect 14924 8032 14976 8041
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 15384 7896 15436 7948
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 12072 7828 12124 7880
rect 14096 7828 14148 7880
rect 14740 7871 14792 7880
rect 14740 7837 14749 7871
rect 14749 7837 14783 7871
rect 14783 7837 14792 7871
rect 14740 7828 14792 7837
rect 14648 7760 14700 7812
rect 11060 7692 11112 7744
rect 13360 7692 13412 7744
rect 13544 7735 13596 7744
rect 13544 7701 13553 7735
rect 13553 7701 13587 7735
rect 13587 7701 13596 7735
rect 13544 7692 13596 7701
rect 6880 7590 6932 7642
rect 6944 7590 6996 7642
rect 7008 7590 7060 7642
rect 7072 7590 7124 7642
rect 7136 7590 7188 7642
rect 12811 7590 12863 7642
rect 12875 7590 12927 7642
rect 12939 7590 12991 7642
rect 13003 7590 13055 7642
rect 13067 7590 13119 7642
rect 8484 7488 8536 7540
rect 11520 7531 11572 7540
rect 11520 7497 11529 7531
rect 11529 7497 11563 7531
rect 11563 7497 11572 7531
rect 11520 7488 11572 7497
rect 8852 7420 8904 7472
rect 13544 7420 13596 7472
rect 8392 7395 8444 7404
rect 8392 7361 8426 7395
rect 8426 7361 8444 7395
rect 8392 7352 8444 7361
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10692 7352 10744 7361
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 12624 7395 12676 7404
rect 12624 7361 12633 7395
rect 12633 7361 12667 7395
rect 12667 7361 12676 7395
rect 12624 7352 12676 7361
rect 11060 7284 11112 7336
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 14004 7327 14056 7336
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 10232 7148 10284 7200
rect 10876 7148 10928 7200
rect 11980 7148 12032 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 16212 7148 16264 7200
rect 3915 7046 3967 7098
rect 3979 7046 4031 7098
rect 4043 7046 4095 7098
rect 4107 7046 4159 7098
rect 4171 7046 4223 7098
rect 9846 7046 9898 7098
rect 9910 7046 9962 7098
rect 9974 7046 10026 7098
rect 10038 7046 10090 7098
rect 10102 7046 10154 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 15904 7046 15956 7098
rect 15968 7046 16020 7098
rect 16032 7046 16084 7098
rect 8392 6944 8444 6996
rect 14740 6876 14792 6928
rect 7472 6740 7524 6792
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8116 6808 8168 6860
rect 8852 6808 8904 6860
rect 9496 6808 9548 6860
rect 11428 6808 11480 6860
rect 14832 6808 14884 6860
rect 15016 6808 15068 6860
rect 8484 6740 8536 6792
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 12440 6740 12492 6792
rect 14004 6740 14056 6792
rect 15108 6740 15160 6792
rect 14372 6672 14424 6724
rect 14924 6672 14976 6724
rect 16764 6672 16816 6724
rect 9772 6604 9824 6656
rect 12440 6604 12492 6656
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 16212 6604 16264 6656
rect 6880 6502 6932 6554
rect 6944 6502 6996 6554
rect 7008 6502 7060 6554
rect 7072 6502 7124 6554
rect 7136 6502 7188 6554
rect 12811 6502 12863 6554
rect 12875 6502 12927 6554
rect 12939 6502 12991 6554
rect 13003 6502 13055 6554
rect 13067 6502 13119 6554
rect 7748 6400 7800 6452
rect 11612 6400 11664 6452
rect 12440 6443 12492 6452
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 12624 6400 12676 6452
rect 14556 6400 14608 6452
rect 15108 6400 15160 6452
rect 6552 6332 6604 6384
rect 5264 6264 5316 6316
rect 6736 6264 6788 6316
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 12164 6264 12216 6316
rect 12624 6264 12676 6316
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 5540 6196 5592 6248
rect 8116 6196 8168 6248
rect 15568 6264 15620 6316
rect 17316 6307 17368 6316
rect 17316 6273 17325 6307
rect 17325 6273 17359 6307
rect 17359 6273 17368 6307
rect 17316 6264 17368 6273
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 12256 6128 12308 6180
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 7472 6060 7524 6112
rect 16948 6060 17000 6112
rect 3915 5958 3967 6010
rect 3979 5958 4031 6010
rect 4043 5958 4095 6010
rect 4107 5958 4159 6010
rect 4171 5958 4223 6010
rect 9846 5958 9898 6010
rect 9910 5958 9962 6010
rect 9974 5958 10026 6010
rect 10038 5958 10090 6010
rect 10102 5958 10154 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 15904 5958 15956 6010
rect 15968 5958 16020 6010
rect 16032 5958 16084 6010
rect 4988 5856 5040 5908
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 11888 5856 11940 5908
rect 12624 5899 12676 5908
rect 12624 5865 12633 5899
rect 12633 5865 12667 5899
rect 12667 5865 12676 5899
rect 12624 5856 12676 5865
rect 15568 5856 15620 5908
rect 16764 5899 16816 5908
rect 16764 5865 16773 5899
rect 16773 5865 16807 5899
rect 16807 5865 16816 5899
rect 16764 5856 16816 5865
rect 17316 5856 17368 5908
rect 6644 5788 6696 5840
rect 9220 5788 9272 5840
rect 4528 5720 4580 5772
rect 7656 5720 7708 5772
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 12440 5763 12492 5772
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 12440 5720 12492 5729
rect 14740 5720 14792 5772
rect 5080 5695 5132 5704
rect 5080 5661 5089 5695
rect 5089 5661 5123 5695
rect 5123 5661 5132 5695
rect 5080 5652 5132 5661
rect 5540 5652 5592 5704
rect 6644 5652 6696 5704
rect 7564 5652 7616 5704
rect 8300 5695 8352 5704
rect 6736 5584 6788 5636
rect 7288 5584 7340 5636
rect 7748 5584 7800 5636
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 9772 5695 9824 5704
rect 9772 5661 9806 5695
rect 9806 5661 9824 5695
rect 9772 5652 9824 5661
rect 11060 5652 11112 5704
rect 12256 5652 12308 5704
rect 13360 5652 13412 5704
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 5540 5516 5592 5568
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 12164 5584 12216 5636
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16948 5695 17000 5704
rect 16212 5652 16264 5661
rect 16948 5661 16957 5695
rect 16957 5661 16991 5695
rect 16991 5661 17000 5695
rect 16948 5652 17000 5661
rect 17868 5652 17920 5704
rect 13360 5516 13412 5568
rect 14280 5516 14332 5568
rect 14924 5516 14976 5568
rect 15568 5516 15620 5568
rect 6880 5414 6932 5466
rect 6944 5414 6996 5466
rect 7008 5414 7060 5466
rect 7072 5414 7124 5466
rect 7136 5414 7188 5466
rect 12811 5414 12863 5466
rect 12875 5414 12927 5466
rect 12939 5414 12991 5466
rect 13003 5414 13055 5466
rect 13067 5414 13119 5466
rect 5080 5312 5132 5364
rect 8300 5312 8352 5364
rect 12164 5355 12216 5364
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 14740 5312 14792 5364
rect 6736 5287 6788 5296
rect 6736 5253 6745 5287
rect 6745 5253 6779 5287
rect 6779 5253 6788 5287
rect 6736 5244 6788 5253
rect 5448 5108 5500 5160
rect 5356 5040 5408 5092
rect 6644 5176 6696 5228
rect 7380 5244 7432 5296
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 8024 5244 8076 5296
rect 7748 5176 7800 5228
rect 8300 5176 8352 5228
rect 10876 5176 10928 5228
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 13452 5176 13504 5228
rect 14004 5219 14056 5228
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 14740 5176 14792 5228
rect 11060 5108 11112 5160
rect 5540 4972 5592 5024
rect 6368 4972 6420 5024
rect 7564 4972 7616 5024
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 9680 4972 9732 5024
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 3915 4870 3967 4922
rect 3979 4870 4031 4922
rect 4043 4870 4095 4922
rect 4107 4870 4159 4922
rect 4171 4870 4223 4922
rect 9846 4870 9898 4922
rect 9910 4870 9962 4922
rect 9974 4870 10026 4922
rect 10038 4870 10090 4922
rect 10102 4870 10154 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 15904 4870 15956 4922
rect 15968 4870 16020 4922
rect 16032 4870 16084 4922
rect 7656 4768 7708 4820
rect 7748 4768 7800 4820
rect 11152 4768 11204 4820
rect 11796 4768 11848 4820
rect 12624 4768 12676 4820
rect 13452 4768 13504 4820
rect 14740 4811 14792 4820
rect 14740 4777 14749 4811
rect 14749 4777 14783 4811
rect 14783 4777 14792 4811
rect 14740 4768 14792 4777
rect 5540 4632 5592 4684
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 6644 4700 6696 4752
rect 7472 4700 7524 4752
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7380 4564 7432 4616
rect 8116 4632 8168 4684
rect 9496 4632 9548 4684
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 8392 4564 8444 4616
rect 9680 4564 9732 4616
rect 11704 4607 11756 4616
rect 11704 4573 11738 4607
rect 11738 4573 11756 4607
rect 11704 4564 11756 4573
rect 13360 4564 13412 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14924 4607 14976 4616
rect 14924 4573 14933 4607
rect 14933 4573 14967 4607
rect 14967 4573 14976 4607
rect 14924 4564 14976 4573
rect 15568 4607 15620 4616
rect 15568 4573 15577 4607
rect 15577 4573 15611 4607
rect 15611 4573 15620 4607
rect 15568 4564 15620 4573
rect 8300 4539 8352 4548
rect 5724 4471 5776 4480
rect 5724 4437 5733 4471
rect 5733 4437 5767 4471
rect 5767 4437 5776 4471
rect 5724 4428 5776 4437
rect 6184 4471 6236 4480
rect 6184 4437 6193 4471
rect 6193 4437 6227 4471
rect 6227 4437 6236 4471
rect 6184 4428 6236 4437
rect 6552 4428 6604 4480
rect 8300 4505 8309 4539
rect 8309 4505 8343 4539
rect 8343 4505 8352 4539
rect 8300 4496 8352 4505
rect 13268 4471 13320 4480
rect 13268 4437 13277 4471
rect 13277 4437 13311 4471
rect 13311 4437 13320 4471
rect 13268 4428 13320 4437
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 6880 4326 6932 4378
rect 6944 4326 6996 4378
rect 7008 4326 7060 4378
rect 7072 4326 7124 4378
rect 7136 4326 7188 4378
rect 12811 4326 12863 4378
rect 12875 4326 12927 4378
rect 12939 4326 12991 4378
rect 13003 4326 13055 4378
rect 13067 4326 13119 4378
rect 6644 4224 6696 4276
rect 8300 4224 8352 4276
rect 10508 4267 10560 4276
rect 10508 4233 10517 4267
rect 10517 4233 10551 4267
rect 10551 4233 10560 4267
rect 10508 4224 10560 4233
rect 5724 4088 5776 4140
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7564 4131 7616 4140
rect 7564 4097 7598 4131
rect 7598 4097 7616 4131
rect 6092 4020 6144 4072
rect 7564 4088 7616 4097
rect 9496 4156 9548 4208
rect 13268 4156 13320 4208
rect 9772 4088 9824 4140
rect 14004 4088 14056 4140
rect 15384 4156 15436 4208
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 15476 4088 15528 4140
rect 13728 3995 13780 4004
rect 13728 3961 13737 3995
rect 13737 3961 13771 3995
rect 13771 3961 13780 3995
rect 13728 3952 13780 3961
rect 12164 3884 12216 3936
rect 16856 3884 16908 3936
rect 3915 3782 3967 3834
rect 3979 3782 4031 3834
rect 4043 3782 4095 3834
rect 4107 3782 4159 3834
rect 4171 3782 4223 3834
rect 9846 3782 9898 3834
rect 9910 3782 9962 3834
rect 9974 3782 10026 3834
rect 10038 3782 10090 3834
rect 10102 3782 10154 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 15904 3782 15956 3834
rect 15968 3782 16020 3834
rect 16032 3782 16084 3834
rect 7472 3723 7524 3732
rect 7472 3689 7481 3723
rect 7481 3689 7515 3723
rect 7515 3689 7524 3723
rect 7472 3680 7524 3689
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 11520 3680 11572 3732
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 12532 3612 12584 3664
rect 11152 3544 11204 3596
rect 6184 3476 6236 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 11060 3519 11112 3528
rect 11060 3485 11069 3519
rect 11069 3485 11103 3519
rect 11103 3485 11112 3519
rect 11060 3476 11112 3485
rect 6880 3238 6932 3290
rect 6944 3238 6996 3290
rect 7008 3238 7060 3290
rect 7072 3238 7124 3290
rect 7136 3238 7188 3290
rect 12811 3238 12863 3290
rect 12875 3238 12927 3290
rect 12939 3238 12991 3290
rect 13003 3238 13055 3290
rect 13067 3238 13119 3290
rect 3915 2694 3967 2746
rect 3979 2694 4031 2746
rect 4043 2694 4095 2746
rect 4107 2694 4159 2746
rect 4171 2694 4223 2746
rect 9846 2694 9898 2746
rect 9910 2694 9962 2746
rect 9974 2694 10026 2746
rect 10038 2694 10090 2746
rect 10102 2694 10154 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 15904 2694 15956 2746
rect 15968 2694 16020 2746
rect 16032 2694 16084 2746
rect 9128 2592 9180 2644
rect 20 2388 72 2440
rect 8392 2388 8444 2440
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 16764 2252 16816 2304
rect 6880 2150 6932 2202
rect 6944 2150 6996 2202
rect 7008 2150 7060 2202
rect 7072 2150 7124 2202
rect 7136 2150 7188 2202
rect 12811 2150 12863 2202
rect 12875 2150 12927 2202
rect 12939 2150 12991 2202
rect 13003 2150 13055 2202
rect 13067 2150 13119 2202
<< metal2 >>
rect 2594 49314 2650 50000
rect 2594 49286 2728 49314
rect 2594 49200 2650 49286
rect 2700 48090 2728 49286
rect 10966 49200 11022 50000
rect 19338 49200 19394 50000
rect 2700 48062 2820 48090
rect 2792 47054 2820 48062
rect 3915 47356 4223 47376
rect 3915 47354 3921 47356
rect 3977 47354 4001 47356
rect 4057 47354 4081 47356
rect 4137 47354 4161 47356
rect 4217 47354 4223 47356
rect 3977 47302 3979 47354
rect 4159 47302 4161 47354
rect 3915 47300 3921 47302
rect 3977 47300 4001 47302
rect 4057 47300 4081 47302
rect 4137 47300 4161 47302
rect 4217 47300 4223 47302
rect 3915 47280 4223 47300
rect 9846 47356 10154 47376
rect 9846 47354 9852 47356
rect 9908 47354 9932 47356
rect 9988 47354 10012 47356
rect 10068 47354 10092 47356
rect 10148 47354 10154 47356
rect 9908 47302 9910 47354
rect 10090 47302 10092 47354
rect 9846 47300 9852 47302
rect 9908 47300 9932 47302
rect 9988 47300 10012 47302
rect 10068 47300 10092 47302
rect 10148 47300 10154 47302
rect 9846 47280 10154 47300
rect 10980 47274 11008 49200
rect 15776 47356 16084 47376
rect 15776 47354 15782 47356
rect 15838 47354 15862 47356
rect 15918 47354 15942 47356
rect 15998 47354 16022 47356
rect 16078 47354 16084 47356
rect 15838 47302 15840 47354
rect 16020 47302 16022 47354
rect 15776 47300 15782 47302
rect 15838 47300 15862 47302
rect 15918 47300 15942 47302
rect 15998 47300 16022 47302
rect 16078 47300 16084 47302
rect 15776 47280 16084 47300
rect 10980 47258 11100 47274
rect 19352 47258 19380 49200
rect 10980 47252 11112 47258
rect 10980 47246 11060 47252
rect 11060 47194 11112 47200
rect 19340 47252 19392 47258
rect 19340 47194 19392 47200
rect 2780 47048 2832 47054
rect 2780 46990 2832 46996
rect 17868 47048 17920 47054
rect 17868 46990 17920 46996
rect 3240 46980 3292 46986
rect 3240 46922 3292 46928
rect 1860 44396 1912 44402
rect 1860 44338 1912 44344
rect 1872 44305 1900 44338
rect 1858 44296 1914 44305
rect 1858 44231 1914 44240
rect 2780 37868 2832 37874
rect 2780 37810 2832 37816
rect 2792 37126 2820 37810
rect 3148 37800 3200 37806
rect 3148 37742 3200 37748
rect 2964 37664 3016 37670
rect 2964 37606 3016 37612
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 2792 36786 2820 37062
rect 2780 36780 2832 36786
rect 2780 36722 2832 36728
rect 2976 36718 3004 37606
rect 3160 37262 3188 37742
rect 3148 37256 3200 37262
rect 3148 37198 3200 37204
rect 2688 36712 2740 36718
rect 2688 36654 2740 36660
rect 2964 36712 3016 36718
rect 2964 36654 3016 36660
rect 1400 35624 1452 35630
rect 1400 35566 1452 35572
rect 1676 35624 1728 35630
rect 1676 35566 1728 35572
rect 1412 35465 1440 35566
rect 1398 35456 1454 35465
rect 1398 35391 1454 35400
rect 1492 26784 1544 26790
rect 1492 26726 1544 26732
rect 1504 26625 1532 26726
rect 1490 26616 1546 26625
rect 1490 26551 1546 26560
rect 1688 26518 1716 35566
rect 2596 31272 2648 31278
rect 2596 31214 2648 31220
rect 2608 29102 2636 31214
rect 2700 30938 2728 36654
rect 3160 36378 3188 37198
rect 3148 36372 3200 36378
rect 3148 36314 3200 36320
rect 3056 31476 3108 31482
rect 3056 31418 3108 31424
rect 2688 30932 2740 30938
rect 2688 30874 2740 30880
rect 3068 30870 3096 31418
rect 3056 30864 3108 30870
rect 3056 30806 3108 30812
rect 2872 30728 2924 30734
rect 2872 30670 2924 30676
rect 2964 30728 3016 30734
rect 2964 30670 3016 30676
rect 2884 29646 2912 30670
rect 2976 29714 3004 30670
rect 2964 29708 3016 29714
rect 2964 29650 3016 29656
rect 2872 29640 2924 29646
rect 2872 29582 2924 29588
rect 2884 29102 2912 29582
rect 2976 29306 3004 29650
rect 2964 29300 3016 29306
rect 2964 29242 3016 29248
rect 2596 29096 2648 29102
rect 2596 29038 2648 29044
rect 2872 29096 2924 29102
rect 2872 29038 2924 29044
rect 2608 28994 2636 29038
rect 2424 28966 2636 28994
rect 1676 26512 1728 26518
rect 1676 26454 1728 26460
rect 2424 24274 2452 28966
rect 3252 25430 3280 46922
rect 6880 46812 7188 46832
rect 6880 46810 6886 46812
rect 6942 46810 6966 46812
rect 7022 46810 7046 46812
rect 7102 46810 7126 46812
rect 7182 46810 7188 46812
rect 6942 46758 6944 46810
rect 7124 46758 7126 46810
rect 6880 46756 6886 46758
rect 6942 46756 6966 46758
rect 7022 46756 7046 46758
rect 7102 46756 7126 46758
rect 7182 46756 7188 46758
rect 6880 46736 7188 46756
rect 12811 46812 13119 46832
rect 12811 46810 12817 46812
rect 12873 46810 12897 46812
rect 12953 46810 12977 46812
rect 13033 46810 13057 46812
rect 13113 46810 13119 46812
rect 12873 46758 12875 46810
rect 13055 46758 13057 46810
rect 12811 46756 12817 46758
rect 12873 46756 12897 46758
rect 12953 46756 12977 46758
rect 13033 46756 13057 46758
rect 13113 46756 13119 46758
rect 12811 46736 13119 46756
rect 3915 46268 4223 46288
rect 3915 46266 3921 46268
rect 3977 46266 4001 46268
rect 4057 46266 4081 46268
rect 4137 46266 4161 46268
rect 4217 46266 4223 46268
rect 3977 46214 3979 46266
rect 4159 46214 4161 46266
rect 3915 46212 3921 46214
rect 3977 46212 4001 46214
rect 4057 46212 4081 46214
rect 4137 46212 4161 46214
rect 4217 46212 4223 46214
rect 3915 46192 4223 46212
rect 9846 46268 10154 46288
rect 9846 46266 9852 46268
rect 9908 46266 9932 46268
rect 9988 46266 10012 46268
rect 10068 46266 10092 46268
rect 10148 46266 10154 46268
rect 9908 46214 9910 46266
rect 10090 46214 10092 46266
rect 9846 46212 9852 46214
rect 9908 46212 9932 46214
rect 9988 46212 10012 46214
rect 10068 46212 10092 46214
rect 10148 46212 10154 46214
rect 9846 46192 10154 46212
rect 15776 46268 16084 46288
rect 15776 46266 15782 46268
rect 15838 46266 15862 46268
rect 15918 46266 15942 46268
rect 15998 46266 16022 46268
rect 16078 46266 16084 46268
rect 15838 46214 15840 46266
rect 16020 46214 16022 46266
rect 15776 46212 15782 46214
rect 15838 46212 15862 46214
rect 15918 46212 15942 46214
rect 15998 46212 16022 46214
rect 16078 46212 16084 46214
rect 15776 46192 16084 46212
rect 8852 45960 8904 45966
rect 8852 45902 8904 45908
rect 9128 45960 9180 45966
rect 9128 45902 9180 45908
rect 6880 45724 7188 45744
rect 6880 45722 6886 45724
rect 6942 45722 6966 45724
rect 7022 45722 7046 45724
rect 7102 45722 7126 45724
rect 7182 45722 7188 45724
rect 6942 45670 6944 45722
rect 7124 45670 7126 45722
rect 6880 45668 6886 45670
rect 6942 45668 6966 45670
rect 7022 45668 7046 45670
rect 7102 45668 7126 45670
rect 7182 45668 7188 45670
rect 6880 45648 7188 45668
rect 8864 45558 8892 45902
rect 8852 45552 8904 45558
rect 8852 45494 8904 45500
rect 6184 45416 6236 45422
rect 6184 45358 6236 45364
rect 7932 45416 7984 45422
rect 7932 45358 7984 45364
rect 8116 45416 8168 45422
rect 8116 45358 8168 45364
rect 3915 45180 4223 45200
rect 3915 45178 3921 45180
rect 3977 45178 4001 45180
rect 4057 45178 4081 45180
rect 4137 45178 4161 45180
rect 4217 45178 4223 45180
rect 3977 45126 3979 45178
rect 4159 45126 4161 45178
rect 3915 45124 3921 45126
rect 3977 45124 4001 45126
rect 4057 45124 4081 45126
rect 4137 45124 4161 45126
rect 4217 45124 4223 45126
rect 3915 45104 4223 45124
rect 5816 44804 5868 44810
rect 5816 44746 5868 44752
rect 5828 44538 5856 44746
rect 5816 44532 5868 44538
rect 5816 44474 5868 44480
rect 5816 44396 5868 44402
rect 5816 44338 5868 44344
rect 3915 44092 4223 44112
rect 3915 44090 3921 44092
rect 3977 44090 4001 44092
rect 4057 44090 4081 44092
rect 4137 44090 4161 44092
rect 4217 44090 4223 44092
rect 3977 44038 3979 44090
rect 4159 44038 4161 44090
rect 3915 44036 3921 44038
rect 3977 44036 4001 44038
rect 4057 44036 4081 44038
rect 4137 44036 4161 44038
rect 4217 44036 4223 44038
rect 3915 44016 4223 44036
rect 5828 43994 5856 44338
rect 5816 43988 5868 43994
rect 5816 43930 5868 43936
rect 6196 43858 6224 45358
rect 6920 45280 6972 45286
rect 6920 45222 6972 45228
rect 7472 45280 7524 45286
rect 7472 45222 7524 45228
rect 6932 45082 6960 45222
rect 6920 45076 6972 45082
rect 6920 45018 6972 45024
rect 7380 45076 7432 45082
rect 7380 45018 7432 45024
rect 6368 44872 6420 44878
rect 6368 44814 6420 44820
rect 6184 43852 6236 43858
rect 6184 43794 6236 43800
rect 3915 43004 4223 43024
rect 3915 43002 3921 43004
rect 3977 43002 4001 43004
rect 4057 43002 4081 43004
rect 4137 43002 4161 43004
rect 4217 43002 4223 43004
rect 3977 42950 3979 43002
rect 4159 42950 4161 43002
rect 3915 42948 3921 42950
rect 3977 42948 4001 42950
rect 4057 42948 4081 42950
rect 4137 42948 4161 42950
rect 4217 42948 4223 42950
rect 3915 42928 4223 42948
rect 6196 42838 6224 43794
rect 6380 43790 6408 44814
rect 6552 44736 6604 44742
rect 6552 44678 6604 44684
rect 6460 43920 6512 43926
rect 6460 43862 6512 43868
rect 6368 43784 6420 43790
rect 6368 43726 6420 43732
rect 6184 42832 6236 42838
rect 6184 42774 6236 42780
rect 3915 41916 4223 41936
rect 3915 41914 3921 41916
rect 3977 41914 4001 41916
rect 4057 41914 4081 41916
rect 4137 41914 4161 41916
rect 4217 41914 4223 41916
rect 3977 41862 3979 41914
rect 4159 41862 4161 41914
rect 3915 41860 3921 41862
rect 3977 41860 4001 41862
rect 4057 41860 4081 41862
rect 4137 41860 4161 41862
rect 4217 41860 4223 41862
rect 3915 41840 4223 41860
rect 3915 40828 4223 40848
rect 3915 40826 3921 40828
rect 3977 40826 4001 40828
rect 4057 40826 4081 40828
rect 4137 40826 4161 40828
rect 4217 40826 4223 40828
rect 3977 40774 3979 40826
rect 4159 40774 4161 40826
rect 3915 40772 3921 40774
rect 3977 40772 4001 40774
rect 4057 40772 4081 40774
rect 4137 40772 4161 40774
rect 4217 40772 4223 40774
rect 3915 40752 4223 40772
rect 5632 40044 5684 40050
rect 5632 39986 5684 39992
rect 5540 39840 5592 39846
rect 5540 39782 5592 39788
rect 3915 39740 4223 39760
rect 3915 39738 3921 39740
rect 3977 39738 4001 39740
rect 4057 39738 4081 39740
rect 4137 39738 4161 39740
rect 4217 39738 4223 39740
rect 3977 39686 3979 39738
rect 4159 39686 4161 39738
rect 3915 39684 3921 39686
rect 3977 39684 4001 39686
rect 4057 39684 4081 39686
rect 4137 39684 4161 39686
rect 4217 39684 4223 39686
rect 3915 39664 4223 39684
rect 3608 39432 3660 39438
rect 3608 39374 3660 39380
rect 3620 38962 3648 39374
rect 3608 38956 3660 38962
rect 3608 38898 3660 38904
rect 3700 38956 3752 38962
rect 3700 38898 3752 38904
rect 3712 37194 3740 38898
rect 4528 38752 4580 38758
rect 4528 38694 4580 38700
rect 3915 38652 4223 38672
rect 3915 38650 3921 38652
rect 3977 38650 4001 38652
rect 4057 38650 4081 38652
rect 4137 38650 4161 38652
rect 4217 38650 4223 38652
rect 3977 38598 3979 38650
rect 4159 38598 4161 38650
rect 3915 38596 3921 38598
rect 3977 38596 4001 38598
rect 4057 38596 4081 38598
rect 4137 38596 4161 38598
rect 4217 38596 4223 38598
rect 3915 38576 4223 38596
rect 3792 38344 3844 38350
rect 3792 38286 3844 38292
rect 3608 37188 3660 37194
rect 3608 37130 3660 37136
rect 3700 37188 3752 37194
rect 3700 37130 3752 37136
rect 3620 36718 3648 37130
rect 3804 36922 3832 38286
rect 4252 38208 4304 38214
rect 4252 38150 4304 38156
rect 3915 37564 4223 37584
rect 3915 37562 3921 37564
rect 3977 37562 4001 37564
rect 4057 37562 4081 37564
rect 4137 37562 4161 37564
rect 4217 37562 4223 37564
rect 3977 37510 3979 37562
rect 4159 37510 4161 37562
rect 3915 37508 3921 37510
rect 3977 37508 4001 37510
rect 4057 37508 4081 37510
rect 4137 37508 4161 37510
rect 4217 37508 4223 37510
rect 3915 37488 4223 37508
rect 4264 37262 4292 38150
rect 4252 37256 4304 37262
rect 4252 37198 4304 37204
rect 4436 37256 4488 37262
rect 4436 37198 4488 37204
rect 3792 36916 3844 36922
rect 3792 36858 3844 36864
rect 3608 36712 3660 36718
rect 3608 36654 3660 36660
rect 3620 36106 3648 36654
rect 3915 36476 4223 36496
rect 3915 36474 3921 36476
rect 3977 36474 4001 36476
rect 4057 36474 4081 36476
rect 4137 36474 4161 36476
rect 4217 36474 4223 36476
rect 3977 36422 3979 36474
rect 4159 36422 4161 36474
rect 3915 36420 3921 36422
rect 3977 36420 4001 36422
rect 4057 36420 4081 36422
rect 4137 36420 4161 36422
rect 4217 36420 4223 36422
rect 3915 36400 4223 36420
rect 3608 36100 3660 36106
rect 3608 36042 3660 36048
rect 3620 31278 3648 36042
rect 3915 35388 4223 35408
rect 3915 35386 3921 35388
rect 3977 35386 4001 35388
rect 4057 35386 4081 35388
rect 4137 35386 4161 35388
rect 4217 35386 4223 35388
rect 3977 35334 3979 35386
rect 4159 35334 4161 35386
rect 3915 35332 3921 35334
rect 3977 35332 4001 35334
rect 4057 35332 4081 35334
rect 4137 35332 4161 35334
rect 4217 35332 4223 35334
rect 3915 35312 4223 35332
rect 4448 34490 4476 37198
rect 4540 37194 4568 38694
rect 4896 38344 4948 38350
rect 4896 38286 4948 38292
rect 4712 37868 4764 37874
rect 4712 37810 4764 37816
rect 4528 37188 4580 37194
rect 4528 37130 4580 37136
rect 4540 36242 4568 37130
rect 4724 36854 4752 37810
rect 4908 37398 4936 38286
rect 5552 38282 5580 39782
rect 5644 38434 5672 39986
rect 6000 39976 6052 39982
rect 6000 39918 6052 39924
rect 5908 39840 5960 39846
rect 5908 39782 5960 39788
rect 5920 39370 5948 39782
rect 5908 39364 5960 39370
rect 5908 39306 5960 39312
rect 5724 39296 5776 39302
rect 5724 39238 5776 39244
rect 5736 38962 5764 39238
rect 6012 38962 6040 39918
rect 6380 39438 6408 43726
rect 6472 43450 6500 43862
rect 6564 43790 6592 44678
rect 6880 44636 7188 44656
rect 6880 44634 6886 44636
rect 6942 44634 6966 44636
rect 7022 44634 7046 44636
rect 7102 44634 7126 44636
rect 7182 44634 7188 44636
rect 6942 44582 6944 44634
rect 7124 44582 7126 44634
rect 6880 44580 6886 44582
rect 6942 44580 6966 44582
rect 7022 44580 7046 44582
rect 7102 44580 7126 44582
rect 7182 44580 7188 44582
rect 6880 44560 7188 44580
rect 7392 44470 7420 45018
rect 7484 44470 7512 45222
rect 7564 44872 7616 44878
rect 7564 44814 7616 44820
rect 7380 44464 7432 44470
rect 7380 44406 7432 44412
rect 7472 44464 7524 44470
rect 7472 44406 7524 44412
rect 7472 44192 7524 44198
rect 7472 44134 7524 44140
rect 7484 43790 7512 44134
rect 7576 43994 7604 44814
rect 7944 44538 7972 45358
rect 8024 44872 8076 44878
rect 8024 44814 8076 44820
rect 7932 44532 7984 44538
rect 7932 44474 7984 44480
rect 7840 44396 7892 44402
rect 7840 44338 7892 44344
rect 7748 44328 7800 44334
rect 7748 44270 7800 44276
rect 7564 43988 7616 43994
rect 7564 43930 7616 43936
rect 7760 43790 7788 44270
rect 6552 43784 6604 43790
rect 6552 43726 6604 43732
rect 7472 43784 7524 43790
rect 7472 43726 7524 43732
rect 7748 43784 7800 43790
rect 7748 43726 7800 43732
rect 6460 43444 6512 43450
rect 6460 43386 6512 43392
rect 6472 40390 6500 43386
rect 6564 43110 6592 43726
rect 6880 43548 7188 43568
rect 6880 43546 6886 43548
rect 6942 43546 6966 43548
rect 7022 43546 7046 43548
rect 7102 43546 7126 43548
rect 7182 43546 7188 43548
rect 6942 43494 6944 43546
rect 7124 43494 7126 43546
rect 6880 43492 6886 43494
rect 6942 43492 6966 43494
rect 7022 43492 7046 43494
rect 7102 43492 7126 43494
rect 7182 43492 7188 43494
rect 6880 43472 7188 43492
rect 6552 43104 6604 43110
rect 6552 43046 6604 43052
rect 7748 43104 7800 43110
rect 7748 43046 7800 43052
rect 6880 42460 7188 42480
rect 6880 42458 6886 42460
rect 6942 42458 6966 42460
rect 7022 42458 7046 42460
rect 7102 42458 7126 42460
rect 7182 42458 7188 42460
rect 6942 42406 6944 42458
rect 7124 42406 7126 42458
rect 6880 42404 6886 42406
rect 6942 42404 6966 42406
rect 7022 42404 7046 42406
rect 7102 42404 7126 42406
rect 7182 42404 7188 42406
rect 6880 42384 7188 42404
rect 7656 42220 7708 42226
rect 7656 42162 7708 42168
rect 6880 41372 7188 41392
rect 6880 41370 6886 41372
rect 6942 41370 6966 41372
rect 7022 41370 7046 41372
rect 7102 41370 7126 41372
rect 7182 41370 7188 41372
rect 6942 41318 6944 41370
rect 7124 41318 7126 41370
rect 6880 41316 6886 41318
rect 6942 41316 6966 41318
rect 7022 41316 7046 41318
rect 7102 41316 7126 41318
rect 7182 41316 7188 41318
rect 6880 41296 7188 41316
rect 6644 40724 6696 40730
rect 6644 40666 6696 40672
rect 6460 40384 6512 40390
rect 6460 40326 6512 40332
rect 6368 39432 6420 39438
rect 6368 39374 6420 39380
rect 6380 39030 6408 39374
rect 6368 39024 6420 39030
rect 6368 38966 6420 38972
rect 5724 38956 5776 38962
rect 5724 38898 5776 38904
rect 6000 38956 6052 38962
rect 6000 38898 6052 38904
rect 6380 38894 6408 38966
rect 6368 38888 6420 38894
rect 6368 38830 6420 38836
rect 5644 38406 5764 38434
rect 5540 38276 5592 38282
rect 5540 38218 5592 38224
rect 5632 38276 5684 38282
rect 5632 38218 5684 38224
rect 5644 37942 5672 38218
rect 5632 37936 5684 37942
rect 5632 37878 5684 37884
rect 5080 37664 5132 37670
rect 5080 37606 5132 37612
rect 5356 37664 5408 37670
rect 5356 37606 5408 37612
rect 4896 37392 4948 37398
rect 4896 37334 4948 37340
rect 4712 36848 4764 36854
rect 4712 36790 4764 36796
rect 4908 36768 4936 37334
rect 4988 37324 5040 37330
rect 4988 37266 5040 37272
rect 5000 36922 5028 37266
rect 5092 37262 5120 37606
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 4988 36916 5040 36922
rect 4988 36858 5040 36864
rect 5368 36786 5396 37606
rect 5736 37194 5764 38406
rect 6380 38350 6408 38830
rect 6368 38344 6420 38350
rect 6368 38286 6420 38292
rect 6472 37194 6500 40326
rect 6656 40050 6684 40666
rect 6736 40452 6788 40458
rect 6736 40394 6788 40400
rect 6552 40044 6604 40050
rect 6552 39986 6604 39992
rect 6644 40044 6696 40050
rect 6644 39986 6696 39992
rect 6564 39098 6592 39986
rect 6748 39982 6776 40394
rect 6880 40284 7188 40304
rect 6880 40282 6886 40284
rect 6942 40282 6966 40284
rect 7022 40282 7046 40284
rect 7102 40282 7126 40284
rect 7182 40282 7188 40284
rect 6942 40230 6944 40282
rect 7124 40230 7126 40282
rect 6880 40228 6886 40230
rect 6942 40228 6966 40230
rect 7022 40228 7046 40230
rect 7102 40228 7126 40230
rect 7182 40228 7188 40230
rect 6880 40208 7188 40228
rect 6736 39976 6788 39982
rect 6736 39918 6788 39924
rect 6828 39976 6880 39982
rect 6828 39918 6880 39924
rect 6840 39370 6868 39918
rect 7564 39568 7616 39574
rect 7564 39510 7616 39516
rect 7380 39500 7432 39506
rect 7380 39442 7432 39448
rect 6828 39364 6880 39370
rect 6828 39306 6880 39312
rect 6880 39196 7188 39216
rect 6880 39194 6886 39196
rect 6942 39194 6966 39196
rect 7022 39194 7046 39196
rect 7102 39194 7126 39196
rect 7182 39194 7188 39196
rect 6942 39142 6944 39194
rect 7124 39142 7126 39194
rect 6880 39140 6886 39142
rect 6942 39140 6966 39142
rect 7022 39140 7046 39142
rect 7102 39140 7126 39142
rect 7182 39140 7188 39142
rect 6880 39120 7188 39140
rect 6552 39092 6604 39098
rect 6552 39034 6604 39040
rect 7288 39024 7340 39030
rect 7288 38966 7340 38972
rect 6644 38956 6696 38962
rect 6644 38898 6696 38904
rect 6552 37868 6604 37874
rect 6552 37810 6604 37816
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5724 37188 5776 37194
rect 5724 37130 5776 37136
rect 6460 37188 6512 37194
rect 6460 37130 6512 37136
rect 5448 37120 5500 37126
rect 5448 37062 5500 37068
rect 5460 36854 5488 37062
rect 5448 36848 5500 36854
rect 5448 36790 5500 36796
rect 5080 36780 5132 36786
rect 4908 36740 5080 36768
rect 5080 36722 5132 36728
rect 5356 36780 5408 36786
rect 5356 36722 5408 36728
rect 4620 36712 4672 36718
rect 4620 36654 4672 36660
rect 4528 36236 4580 36242
rect 4528 36178 4580 36184
rect 4540 35698 4568 36178
rect 4528 35692 4580 35698
rect 4528 35634 4580 35640
rect 4356 34462 4476 34490
rect 3915 34300 4223 34320
rect 3915 34298 3921 34300
rect 3977 34298 4001 34300
rect 4057 34298 4081 34300
rect 4137 34298 4161 34300
rect 4217 34298 4223 34300
rect 3977 34246 3979 34298
rect 4159 34246 4161 34298
rect 3915 34244 3921 34246
rect 3977 34244 4001 34246
rect 4057 34244 4081 34246
rect 4137 34244 4161 34246
rect 4217 34244 4223 34246
rect 3915 34224 4223 34244
rect 3915 33212 4223 33232
rect 3915 33210 3921 33212
rect 3977 33210 4001 33212
rect 4057 33210 4081 33212
rect 4137 33210 4161 33212
rect 4217 33210 4223 33212
rect 3977 33158 3979 33210
rect 4159 33158 4161 33210
rect 3915 33156 3921 33158
rect 3977 33156 4001 33158
rect 4057 33156 4081 33158
rect 4137 33156 4161 33158
rect 4217 33156 4223 33158
rect 3915 33136 4223 33156
rect 3700 32904 3752 32910
rect 3700 32846 3752 32852
rect 3608 31272 3660 31278
rect 3608 31214 3660 31220
rect 3516 31136 3568 31142
rect 3516 31078 3568 31084
rect 3528 30734 3556 31078
rect 3620 30734 3648 31214
rect 3516 30728 3568 30734
rect 3516 30670 3568 30676
rect 3608 30728 3660 30734
rect 3608 30670 3660 30676
rect 3332 29096 3384 29102
rect 3332 29038 3384 29044
rect 3240 25424 3292 25430
rect 3240 25366 3292 25372
rect 2412 24268 2464 24274
rect 2412 24210 2464 24216
rect 2964 24064 3016 24070
rect 2964 24006 3016 24012
rect 3148 24064 3200 24070
rect 3148 24006 3200 24012
rect 2976 23730 3004 24006
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 2976 23254 3004 23666
rect 2964 23248 3016 23254
rect 2964 23190 3016 23196
rect 3160 23118 3188 24006
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 3252 23186 3280 23666
rect 3344 23322 3372 29038
rect 3608 28552 3660 28558
rect 3608 28494 3660 28500
rect 3620 26450 3648 28494
rect 3608 26444 3660 26450
rect 3608 26386 3660 26392
rect 3620 25906 3648 26386
rect 3712 26234 3740 32846
rect 4252 32836 4304 32842
rect 4252 32778 4304 32784
rect 3884 32768 3936 32774
rect 3884 32710 3936 32716
rect 3896 32434 3924 32710
rect 3884 32428 3936 32434
rect 3884 32370 3936 32376
rect 3915 32124 4223 32144
rect 3915 32122 3921 32124
rect 3977 32122 4001 32124
rect 4057 32122 4081 32124
rect 4137 32122 4161 32124
rect 4217 32122 4223 32124
rect 3977 32070 3979 32122
rect 4159 32070 4161 32122
rect 3915 32068 3921 32070
rect 3977 32068 4001 32070
rect 4057 32068 4081 32070
rect 4137 32068 4161 32070
rect 4217 32068 4223 32070
rect 3915 32048 4223 32068
rect 4264 32026 4292 32778
rect 4252 32020 4304 32026
rect 4252 31962 4304 31968
rect 3792 31884 3844 31890
rect 3792 31826 3844 31832
rect 3804 30938 3832 31826
rect 3976 31816 4028 31822
rect 3976 31758 4028 31764
rect 3988 31482 4016 31758
rect 3976 31476 4028 31482
rect 3976 31418 4028 31424
rect 4252 31136 4304 31142
rect 4252 31078 4304 31084
rect 3915 31036 4223 31056
rect 3915 31034 3921 31036
rect 3977 31034 4001 31036
rect 4057 31034 4081 31036
rect 4137 31034 4161 31036
rect 4217 31034 4223 31036
rect 3977 30982 3979 31034
rect 4159 30982 4161 31034
rect 3915 30980 3921 30982
rect 3977 30980 4001 30982
rect 4057 30980 4081 30982
rect 4137 30980 4161 30982
rect 4217 30980 4223 30982
rect 3915 30960 4223 30980
rect 3792 30932 3844 30938
rect 3792 30874 3844 30880
rect 4264 30598 4292 31078
rect 3792 30592 3844 30598
rect 3792 30534 3844 30540
rect 4252 30592 4304 30598
rect 4252 30534 4304 30540
rect 3804 29782 3832 30534
rect 3915 29948 4223 29968
rect 3915 29946 3921 29948
rect 3977 29946 4001 29948
rect 4057 29946 4081 29948
rect 4137 29946 4161 29948
rect 4217 29946 4223 29948
rect 3977 29894 3979 29946
rect 4159 29894 4161 29946
rect 3915 29892 3921 29894
rect 3977 29892 4001 29894
rect 4057 29892 4081 29894
rect 4137 29892 4161 29894
rect 4217 29892 4223 29894
rect 3915 29872 4223 29892
rect 3792 29776 3844 29782
rect 4264 29730 4292 30534
rect 3792 29718 3844 29724
rect 3804 29170 3832 29718
rect 4172 29702 4292 29730
rect 3792 29164 3844 29170
rect 3792 29106 3844 29112
rect 4172 29034 4200 29702
rect 4160 29028 4212 29034
rect 4160 28970 4212 28976
rect 4356 28994 4384 34462
rect 4436 33312 4488 33318
rect 4436 33254 4488 33260
rect 4448 32502 4476 33254
rect 4632 32978 4660 36654
rect 4896 36576 4948 36582
rect 4896 36518 4948 36524
rect 4908 36378 4936 36518
rect 4896 36372 4948 36378
rect 4896 36314 4948 36320
rect 4804 36100 4856 36106
rect 4804 36042 4856 36048
rect 4712 33108 4764 33114
rect 4712 33050 4764 33056
rect 4620 32972 4672 32978
rect 4620 32914 4672 32920
rect 4724 32910 4752 33050
rect 4528 32904 4580 32910
rect 4528 32846 4580 32852
rect 4712 32904 4764 32910
rect 4712 32846 4764 32852
rect 4436 32496 4488 32502
rect 4436 32438 4488 32444
rect 4540 32026 4568 32846
rect 4620 32768 4672 32774
rect 4620 32710 4672 32716
rect 4528 32020 4580 32026
rect 4528 31962 4580 31968
rect 4632 28994 4660 32710
rect 4356 28966 4476 28994
rect 4252 28960 4304 28966
rect 4252 28902 4304 28908
rect 3915 28860 4223 28880
rect 3915 28858 3921 28860
rect 3977 28858 4001 28860
rect 4057 28858 4081 28860
rect 4137 28858 4161 28860
rect 4217 28858 4223 28860
rect 3977 28806 3979 28858
rect 4159 28806 4161 28858
rect 3915 28804 3921 28806
rect 3977 28804 4001 28806
rect 4057 28804 4081 28806
rect 4137 28804 4161 28806
rect 4217 28804 4223 28806
rect 3915 28784 4223 28804
rect 3792 28484 3844 28490
rect 3792 28426 3844 28432
rect 3804 28218 3832 28426
rect 3792 28212 3844 28218
rect 3792 28154 3844 28160
rect 4264 28082 4292 28902
rect 4448 28082 4476 28966
rect 4540 28966 4660 28994
rect 4252 28076 4304 28082
rect 4252 28018 4304 28024
rect 4436 28076 4488 28082
rect 4436 28018 4488 28024
rect 3915 27772 4223 27792
rect 3915 27770 3921 27772
rect 3977 27770 4001 27772
rect 4057 27770 4081 27772
rect 4137 27770 4161 27772
rect 4217 27770 4223 27772
rect 3977 27718 3979 27770
rect 4159 27718 4161 27770
rect 3915 27716 3921 27718
rect 3977 27716 4001 27718
rect 4057 27716 4081 27718
rect 4137 27716 4161 27718
rect 4217 27716 4223 27718
rect 3915 27696 4223 27716
rect 4436 27396 4488 27402
rect 4436 27338 4488 27344
rect 4448 26790 4476 27338
rect 4540 26994 4568 28966
rect 4620 28008 4672 28014
rect 4620 27950 4672 27956
rect 4528 26988 4580 26994
rect 4528 26930 4580 26936
rect 4436 26784 4488 26790
rect 4436 26726 4488 26732
rect 3915 26684 4223 26704
rect 3915 26682 3921 26684
rect 3977 26682 4001 26684
rect 4057 26682 4081 26684
rect 4137 26682 4161 26684
rect 4217 26682 4223 26684
rect 3977 26630 3979 26682
rect 4159 26630 4161 26682
rect 3915 26628 3921 26630
rect 3977 26628 4001 26630
rect 4057 26628 4081 26630
rect 4137 26628 4161 26630
rect 4217 26628 4223 26630
rect 3915 26608 4223 26628
rect 4448 26382 4476 26726
rect 4436 26376 4488 26382
rect 4436 26318 4488 26324
rect 3712 26206 3832 26234
rect 3608 25900 3660 25906
rect 3608 25842 3660 25848
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3712 25498 3740 25842
rect 3700 25492 3752 25498
rect 3700 25434 3752 25440
rect 3700 25288 3752 25294
rect 3700 25230 3752 25236
rect 3712 24138 3740 25230
rect 3700 24132 3752 24138
rect 3700 24074 3752 24080
rect 3700 23724 3752 23730
rect 3700 23666 3752 23672
rect 3424 23520 3476 23526
rect 3424 23462 3476 23468
rect 3436 23322 3464 23462
rect 3332 23316 3384 23322
rect 3332 23258 3384 23264
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 3240 23180 3292 23186
rect 3240 23122 3292 23128
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 2884 22642 2912 23054
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2976 22506 3004 23054
rect 3252 22778 3280 23122
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3332 22636 3384 22642
rect 3332 22578 3384 22584
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 2964 22500 3016 22506
rect 2964 22442 3016 22448
rect 2780 22228 2832 22234
rect 2780 22170 2832 22176
rect 2792 22030 2820 22170
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2976 21894 3004 22442
rect 3252 22234 3280 22510
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 2792 21486 2820 21830
rect 3344 21554 3372 22578
rect 3712 22030 3740 23666
rect 3804 22778 3832 26206
rect 3915 25596 4223 25616
rect 3915 25594 3921 25596
rect 3977 25594 4001 25596
rect 4057 25594 4081 25596
rect 4137 25594 4161 25596
rect 4217 25594 4223 25596
rect 3977 25542 3979 25594
rect 4159 25542 4161 25594
rect 3915 25540 3921 25542
rect 3977 25540 4001 25542
rect 4057 25540 4081 25542
rect 4137 25540 4161 25542
rect 4217 25540 4223 25542
rect 3915 25520 4223 25540
rect 4252 25288 4304 25294
rect 4252 25230 4304 25236
rect 3915 24508 4223 24528
rect 3915 24506 3921 24508
rect 3977 24506 4001 24508
rect 4057 24506 4081 24508
rect 4137 24506 4161 24508
rect 4217 24506 4223 24508
rect 3977 24454 3979 24506
rect 4159 24454 4161 24506
rect 3915 24452 3921 24454
rect 3977 24452 4001 24454
rect 4057 24452 4081 24454
rect 4137 24452 4161 24454
rect 4217 24452 4223 24454
rect 3915 24432 4223 24452
rect 3884 24268 3936 24274
rect 3884 24210 3936 24216
rect 3896 23798 3924 24210
rect 4264 23866 4292 25230
rect 4632 25226 4660 27950
rect 4724 27334 4752 32846
rect 4816 31822 4844 36042
rect 5092 33046 5120 36722
rect 5368 36174 5396 36722
rect 5356 36168 5408 36174
rect 5356 36110 5408 36116
rect 5080 33040 5132 33046
rect 5080 32982 5132 32988
rect 5080 32904 5132 32910
rect 5080 32846 5132 32852
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 5000 31822 5028 32166
rect 5092 32026 5120 32846
rect 5080 32020 5132 32026
rect 5080 31962 5132 31968
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 4816 29102 4844 31758
rect 5000 31346 5028 31758
rect 5448 31748 5500 31754
rect 5448 31690 5500 31696
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 5460 29850 5488 31690
rect 5448 29844 5500 29850
rect 5448 29786 5500 29792
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4816 28994 4844 29038
rect 5264 29028 5316 29034
rect 4816 28966 4936 28994
rect 5264 28970 5316 28976
rect 5552 28994 5580 37130
rect 6564 36922 6592 37810
rect 6656 37466 6684 38898
rect 6736 38480 6788 38486
rect 6736 38422 6788 38428
rect 6748 37942 6776 38422
rect 6880 38108 7188 38128
rect 6880 38106 6886 38108
rect 6942 38106 6966 38108
rect 7022 38106 7046 38108
rect 7102 38106 7126 38108
rect 7182 38106 7188 38108
rect 6942 38054 6944 38106
rect 7124 38054 7126 38106
rect 6880 38052 6886 38054
rect 6942 38052 6966 38054
rect 7022 38052 7046 38054
rect 7102 38052 7126 38054
rect 7182 38052 7188 38054
rect 6880 38032 7188 38052
rect 6736 37936 6788 37942
rect 6736 37878 6788 37884
rect 7300 37466 7328 38966
rect 7392 37874 7420 39442
rect 7380 37868 7432 37874
rect 7380 37810 7432 37816
rect 6644 37460 6696 37466
rect 6644 37402 6696 37408
rect 7288 37460 7340 37466
rect 7288 37402 7340 37408
rect 7300 37346 7328 37402
rect 7576 37398 7604 39510
rect 7564 37392 7616 37398
rect 7300 37318 7420 37346
rect 7564 37334 7616 37340
rect 7288 37188 7340 37194
rect 7288 37130 7340 37136
rect 6880 37020 7188 37040
rect 6880 37018 6886 37020
rect 6942 37018 6966 37020
rect 7022 37018 7046 37020
rect 7102 37018 7126 37020
rect 7182 37018 7188 37020
rect 6942 36966 6944 37018
rect 7124 36966 7126 37018
rect 6880 36964 6886 36966
rect 6942 36964 6966 36966
rect 7022 36964 7046 36966
rect 7102 36964 7126 36966
rect 7182 36964 7188 36966
rect 6880 36944 7188 36964
rect 6552 36916 6604 36922
rect 6552 36858 6604 36864
rect 5632 36644 5684 36650
rect 5632 36586 5684 36592
rect 5644 32978 5672 36586
rect 6880 35932 7188 35952
rect 6880 35930 6886 35932
rect 6942 35930 6966 35932
rect 7022 35930 7046 35932
rect 7102 35930 7126 35932
rect 7182 35930 7188 35932
rect 6942 35878 6944 35930
rect 7124 35878 7126 35930
rect 6880 35876 6886 35878
rect 6942 35876 6966 35878
rect 7022 35876 7046 35878
rect 7102 35876 7126 35878
rect 7182 35876 7188 35878
rect 6880 35856 7188 35876
rect 5724 35488 5776 35494
rect 5724 35430 5776 35436
rect 5632 32972 5684 32978
rect 5632 32914 5684 32920
rect 5644 31822 5672 32914
rect 5736 31822 5764 35430
rect 7300 35222 7328 37130
rect 7392 36854 7420 37318
rect 7472 37324 7524 37330
rect 7472 37266 7524 37272
rect 7484 36922 7512 37266
rect 7564 37188 7616 37194
rect 7564 37130 7616 37136
rect 7472 36916 7524 36922
rect 7472 36858 7524 36864
rect 7380 36848 7432 36854
rect 7576 36802 7604 37130
rect 7380 36790 7432 36796
rect 7484 36774 7604 36802
rect 7288 35216 7340 35222
rect 7288 35158 7340 35164
rect 6880 34844 7188 34864
rect 6880 34842 6886 34844
rect 6942 34842 6966 34844
rect 7022 34842 7046 34844
rect 7102 34842 7126 34844
rect 7182 34842 7188 34844
rect 6942 34790 6944 34842
rect 7124 34790 7126 34842
rect 6880 34788 6886 34790
rect 6942 34788 6966 34790
rect 7022 34788 7046 34790
rect 7102 34788 7126 34790
rect 7182 34788 7188 34790
rect 6880 34768 7188 34788
rect 5908 33992 5960 33998
rect 5828 33940 5908 33946
rect 5828 33934 5960 33940
rect 6460 33992 6512 33998
rect 6460 33934 6512 33940
rect 5828 33918 5948 33934
rect 5828 33454 5856 33918
rect 5908 33856 5960 33862
rect 5908 33798 5960 33804
rect 5920 33590 5948 33798
rect 5908 33584 5960 33590
rect 5908 33526 5960 33532
rect 5816 33448 5868 33454
rect 5816 33390 5868 33396
rect 5828 33318 5856 33390
rect 6472 33318 6500 33934
rect 6644 33856 6696 33862
rect 6644 33798 6696 33804
rect 5816 33312 5868 33318
rect 5816 33254 5868 33260
rect 6460 33312 6512 33318
rect 6460 33254 6512 33260
rect 5828 32910 5856 33254
rect 5998 33144 6054 33153
rect 5998 33079 6054 33088
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 5828 31890 5856 32846
rect 6012 32502 6040 33079
rect 6184 32768 6236 32774
rect 6184 32710 6236 32716
rect 6000 32496 6052 32502
rect 6000 32438 6052 32444
rect 6092 32496 6144 32502
rect 6092 32438 6144 32444
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5632 31816 5684 31822
rect 5632 31758 5684 31764
rect 5724 31816 5776 31822
rect 5724 31758 5776 31764
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5644 29646 5672 31418
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5908 29640 5960 29646
rect 5908 29582 5960 29588
rect 5920 29306 5948 29582
rect 5908 29300 5960 29306
rect 5908 29242 5960 29248
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 4712 27124 4764 27130
rect 4712 27066 4764 27072
rect 4724 26382 4752 27066
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4816 25294 4844 28018
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 4620 25220 4672 25226
rect 4620 25162 4672 25168
rect 4344 24268 4396 24274
rect 4344 24210 4396 24216
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 3884 23792 3936 23798
rect 3884 23734 3936 23740
rect 3915 23420 4223 23440
rect 3915 23418 3921 23420
rect 3977 23418 4001 23420
rect 4057 23418 4081 23420
rect 4137 23418 4161 23420
rect 4217 23418 4223 23420
rect 3977 23366 3979 23418
rect 4159 23366 4161 23418
rect 3915 23364 3921 23366
rect 3977 23364 4001 23366
rect 4057 23364 4081 23366
rect 4137 23364 4161 23366
rect 4217 23364 4223 23366
rect 3915 23344 4223 23364
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 3700 22024 3752 22030
rect 3700 21966 3752 21972
rect 3712 21894 3740 21966
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3804 21570 3832 22714
rect 3915 22332 4223 22352
rect 3915 22330 3921 22332
rect 3977 22330 4001 22332
rect 4057 22330 4081 22332
rect 4137 22330 4161 22332
rect 4217 22330 4223 22332
rect 3977 22278 3979 22330
rect 4159 22278 4161 22330
rect 3915 22276 3921 22278
rect 3977 22276 4001 22278
rect 4057 22276 4081 22278
rect 4137 22276 4161 22278
rect 4217 22276 4223 22278
rect 3915 22256 4223 22276
rect 4356 22030 4384 24210
rect 4436 22636 4488 22642
rect 4436 22578 4488 22584
rect 4344 22024 4396 22030
rect 4344 21966 4396 21972
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3620 21542 3832 21570
rect 4252 21548 4304 21554
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 17785 1440 18022
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 2976 16250 3004 21490
rect 3620 20534 3648 21542
rect 4252 21490 4304 21496
rect 3700 21412 3752 21418
rect 3700 21354 3752 21360
rect 3608 20528 3660 20534
rect 3608 20470 3660 20476
rect 3712 20466 3740 21354
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3804 20874 3832 21286
rect 3915 21244 4223 21264
rect 3915 21242 3921 21244
rect 3977 21242 4001 21244
rect 4057 21242 4081 21244
rect 4137 21242 4161 21244
rect 4217 21242 4223 21244
rect 3977 21190 3979 21242
rect 4159 21190 4161 21242
rect 3915 21188 3921 21190
rect 3977 21188 4001 21190
rect 4057 21188 4081 21190
rect 4137 21188 4161 21190
rect 4217 21188 4223 21190
rect 3915 21168 4223 21188
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 4264 20602 4292 21490
rect 4356 20754 4384 21830
rect 4448 20942 4476 22578
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4540 21486 4568 21966
rect 4632 21690 4660 25162
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 22778 4752 22918
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4528 21480 4580 21486
rect 4528 21422 4580 21428
rect 4540 21146 4568 21422
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4356 20726 4476 20754
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3915 20156 4223 20176
rect 3915 20154 3921 20156
rect 3977 20154 4001 20156
rect 4057 20154 4081 20156
rect 4137 20154 4161 20156
rect 4217 20154 4223 20156
rect 3977 20102 3979 20154
rect 4159 20102 4161 20154
rect 3915 20100 3921 20102
rect 3977 20100 4001 20102
rect 4057 20100 4081 20102
rect 4137 20100 4161 20102
rect 4217 20100 4223 20102
rect 3915 20080 4223 20100
rect 3915 19068 4223 19088
rect 3915 19066 3921 19068
rect 3977 19066 4001 19068
rect 4057 19066 4081 19068
rect 4137 19066 4161 19068
rect 4217 19066 4223 19068
rect 3977 19014 3979 19066
rect 4159 19014 4161 19066
rect 3915 19012 3921 19014
rect 3977 19012 4001 19014
rect 4057 19012 4081 19014
rect 4137 19012 4161 19014
rect 4217 19012 4223 19014
rect 3915 18992 4223 19012
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 3915 17980 4223 18000
rect 3915 17978 3921 17980
rect 3977 17978 4001 17980
rect 4057 17978 4081 17980
rect 4137 17978 4161 17980
rect 4217 17978 4223 17980
rect 3977 17926 3979 17978
rect 4159 17926 4161 17978
rect 3915 17924 3921 17926
rect 3977 17924 4001 17926
rect 4057 17924 4081 17926
rect 4137 17924 4161 17926
rect 4217 17924 4223 17926
rect 3915 17904 4223 17924
rect 4264 17218 4292 18226
rect 4172 17202 4292 17218
rect 4160 17196 4292 17202
rect 4212 17190 4292 17196
rect 4160 17138 4212 17144
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2792 15502 2820 16118
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 3068 15366 3096 15982
rect 3252 15434 3280 16050
rect 3344 15978 3372 16458
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3332 15632 3384 15638
rect 3332 15574 3384 15580
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 3068 14618 3096 15302
rect 3344 15026 3372 15574
rect 3436 15026 3464 15846
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3528 14958 3556 16526
rect 3620 15162 3648 17070
rect 3792 17060 3844 17066
rect 3792 17002 3844 17008
rect 3804 16590 3832 17002
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 3915 16892 4223 16912
rect 3915 16890 3921 16892
rect 3977 16890 4001 16892
rect 4057 16890 4081 16892
rect 4137 16890 4161 16892
rect 4217 16890 4223 16892
rect 3977 16838 3979 16890
rect 4159 16838 4161 16890
rect 3915 16836 3921 16838
rect 3977 16836 4001 16838
rect 4057 16836 4081 16838
rect 4137 16836 4161 16838
rect 4217 16836 4223 16838
rect 3915 16816 4223 16836
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3712 15502 3740 15982
rect 3804 15570 3832 16526
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4172 16114 4200 16390
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 3915 15804 4223 15824
rect 3915 15802 3921 15804
rect 3977 15802 4001 15804
rect 4057 15802 4081 15804
rect 4137 15802 4161 15804
rect 4217 15802 4223 15804
rect 3977 15750 3979 15802
rect 4159 15750 4161 15802
rect 3915 15748 3921 15750
rect 3977 15748 4001 15750
rect 4057 15748 4081 15750
rect 4137 15748 4161 15750
rect 4217 15748 4223 15750
rect 3915 15728 4223 15748
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3712 15162 3740 15438
rect 4264 15434 4292 16934
rect 4356 16590 4384 16934
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3915 14716 4223 14736
rect 3915 14714 3921 14716
rect 3977 14714 4001 14716
rect 4057 14714 4081 14716
rect 4137 14714 4161 14716
rect 4217 14714 4223 14716
rect 3977 14662 3979 14714
rect 4159 14662 4161 14714
rect 3915 14660 3921 14662
rect 3977 14660 4001 14662
rect 4057 14660 4081 14662
rect 4137 14660 4161 14662
rect 4217 14660 4223 14662
rect 3915 14640 4223 14660
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 4264 14414 4292 15030
rect 4448 15026 4476 20726
rect 4632 17814 4660 21626
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 4632 17338 4660 17750
rect 4724 17678 4752 22714
rect 4816 21622 4844 25230
rect 4804 21616 4856 21622
rect 4804 21558 4856 21564
rect 4908 17882 4936 28966
rect 5276 28422 5304 28970
rect 5552 28966 5672 28994
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 5276 28150 5304 28358
rect 5264 28144 5316 28150
rect 5264 28086 5316 28092
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 4988 26988 5040 26994
rect 4988 26930 5040 26936
rect 5000 25702 5028 26930
rect 5080 26376 5132 26382
rect 5080 26318 5132 26324
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 5000 25362 5028 25638
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 5092 24818 5120 26318
rect 5172 26308 5224 26314
rect 5172 26250 5224 26256
rect 5184 24818 5212 26250
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5264 25764 5316 25770
rect 5264 25706 5316 25712
rect 5276 25498 5304 25706
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5368 25294 5396 26182
rect 5356 25288 5408 25294
rect 5356 25230 5408 25236
rect 5368 24818 5396 25230
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5184 24410 5212 24754
rect 5172 24404 5224 24410
rect 5172 24346 5224 24352
rect 5172 22976 5224 22982
rect 5172 22918 5224 22924
rect 5184 22642 5212 22918
rect 5460 22778 5488 27270
rect 5552 26586 5580 28494
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5644 25974 5672 28966
rect 5920 28626 5948 29242
rect 5908 28620 5960 28626
rect 5908 28562 5960 28568
rect 5908 28484 5960 28490
rect 5908 28426 5960 28432
rect 5920 27674 5948 28426
rect 5908 27668 5960 27674
rect 5908 27610 5960 27616
rect 5724 27396 5776 27402
rect 5724 27338 5776 27344
rect 5736 27130 5764 27338
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 6012 26234 6040 32438
rect 6104 31822 6132 32438
rect 6092 31816 6144 31822
rect 6092 31758 6144 31764
rect 6092 29640 6144 29646
rect 6092 29582 6144 29588
rect 6104 28558 6132 29582
rect 6092 28552 6144 28558
rect 6092 28494 6144 28500
rect 6104 28014 6132 28494
rect 6092 28008 6144 28014
rect 6092 27950 6144 27956
rect 5920 26206 6040 26234
rect 5632 25968 5684 25974
rect 5632 25910 5684 25916
rect 5632 25492 5684 25498
rect 5632 25434 5684 25440
rect 5644 25158 5672 25434
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5644 24818 5672 25094
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5540 24744 5592 24750
rect 5540 24686 5592 24692
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5552 21554 5580 24686
rect 5644 23118 5672 24754
rect 5736 23322 5764 25230
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5724 23316 5776 23322
rect 5724 23258 5776 23264
rect 5632 23112 5684 23118
rect 5632 23054 5684 23060
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5736 22098 5764 22374
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5552 18426 5580 21490
rect 5644 21434 5672 21830
rect 5736 21554 5764 22034
rect 5828 21690 5856 24754
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5644 21406 5764 21434
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5644 18970 5672 21286
rect 5736 20466 5764 21406
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4632 17134 4660 17274
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4908 16522 4936 17818
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 17338 5212 17614
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5184 16794 5212 17138
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 5276 15706 5304 18226
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17270 5580 18022
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5460 16114 5488 17070
rect 5736 16454 5764 18702
rect 5828 18086 5856 21490
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5920 17814 5948 26206
rect 6092 23044 6144 23050
rect 6196 23032 6224 32710
rect 6472 32570 6500 33254
rect 6656 32842 6684 33798
rect 6880 33756 7188 33776
rect 6880 33754 6886 33756
rect 6942 33754 6966 33756
rect 7022 33754 7046 33756
rect 7102 33754 7126 33756
rect 7182 33754 7188 33756
rect 6942 33702 6944 33754
rect 7124 33702 7126 33754
rect 6880 33700 6886 33702
rect 6942 33700 6966 33702
rect 7022 33700 7046 33702
rect 7102 33700 7126 33702
rect 7182 33700 7188 33702
rect 6880 33680 7188 33700
rect 7300 33590 7328 35158
rect 7484 33930 7512 36774
rect 7564 33992 7616 33998
rect 7564 33934 7616 33940
rect 7472 33924 7524 33930
rect 7472 33866 7524 33872
rect 7288 33584 7340 33590
rect 7288 33526 7340 33532
rect 7380 33380 7432 33386
rect 7380 33322 7432 33328
rect 7392 32910 7420 33322
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 6644 32836 6696 32842
rect 6644 32778 6696 32784
rect 7288 32768 7340 32774
rect 7288 32710 7340 32716
rect 6880 32668 7188 32688
rect 6880 32666 6886 32668
rect 6942 32666 6966 32668
rect 7022 32666 7046 32668
rect 7102 32666 7126 32668
rect 7182 32666 7188 32668
rect 6942 32614 6944 32666
rect 7124 32614 7126 32666
rect 6880 32612 6886 32614
rect 6942 32612 6966 32614
rect 7022 32612 7046 32614
rect 7102 32612 7126 32614
rect 7182 32612 7188 32614
rect 6880 32592 7188 32612
rect 6460 32564 6512 32570
rect 6460 32506 6512 32512
rect 7104 32496 7156 32502
rect 7104 32438 7156 32444
rect 6920 32224 6972 32230
rect 6920 32166 6972 32172
rect 6736 31816 6788 31822
rect 6736 31758 6788 31764
rect 6748 31482 6776 31758
rect 6932 31754 6960 32166
rect 7012 31952 7064 31958
rect 7012 31894 7064 31900
rect 7024 31822 7052 31894
rect 7116 31822 7144 32438
rect 7300 32434 7328 32710
rect 7288 32428 7340 32434
rect 7288 32370 7340 32376
rect 7288 32292 7340 32298
rect 7288 32234 7340 32240
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 6920 31748 6972 31754
rect 6920 31690 6972 31696
rect 6880 31580 7188 31600
rect 6880 31578 6886 31580
rect 6942 31578 6966 31580
rect 7022 31578 7046 31580
rect 7102 31578 7126 31580
rect 7182 31578 7188 31580
rect 6942 31526 6944 31578
rect 7124 31526 7126 31578
rect 6880 31524 6886 31526
rect 6942 31524 6966 31526
rect 7022 31524 7046 31526
rect 7102 31524 7126 31526
rect 7182 31524 7188 31526
rect 6880 31504 7188 31524
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 7300 31414 7328 32234
rect 7288 31408 7340 31414
rect 7288 31350 7340 31356
rect 6828 31136 6880 31142
rect 6828 31078 6880 31084
rect 7196 31136 7248 31142
rect 7196 31078 7248 31084
rect 6840 30666 6868 31078
rect 7208 30666 7236 31078
rect 7392 30818 7420 32846
rect 7576 32570 7604 33934
rect 7564 32564 7616 32570
rect 7564 32506 7616 32512
rect 7472 32360 7524 32366
rect 7472 32302 7524 32308
rect 7484 32026 7512 32302
rect 7472 32020 7524 32026
rect 7472 31962 7524 31968
rect 7668 31754 7696 42162
rect 7760 40526 7788 43046
rect 7852 42226 7880 44338
rect 7944 43382 7972 44474
rect 7932 43376 7984 43382
rect 7932 43318 7984 43324
rect 8036 43194 8064 44814
rect 8128 44266 8156 45358
rect 8864 45354 8892 45494
rect 8852 45348 8904 45354
rect 8852 45290 8904 45296
rect 8668 45280 8720 45286
rect 8668 45222 8720 45228
rect 9036 45280 9088 45286
rect 9036 45222 9088 45228
rect 8300 44872 8352 44878
rect 8300 44814 8352 44820
rect 8116 44260 8168 44266
rect 8116 44202 8168 44208
rect 8128 43314 8156 44202
rect 8116 43308 8168 43314
rect 8116 43250 8168 43256
rect 7944 43166 8064 43194
rect 7840 42220 7892 42226
rect 7840 42162 7892 42168
rect 7944 42022 7972 43166
rect 8312 43110 8340 44814
rect 8392 44736 8444 44742
rect 8392 44678 8444 44684
rect 8404 44402 8432 44678
rect 8680 44402 8708 45222
rect 9048 44878 9076 45222
rect 8944 44872 8996 44878
rect 8944 44814 8996 44820
rect 9036 44872 9088 44878
rect 9036 44814 9088 44820
rect 8392 44396 8444 44402
rect 8392 44338 8444 44344
rect 8668 44396 8720 44402
rect 8668 44338 8720 44344
rect 8680 43994 8708 44338
rect 8668 43988 8720 43994
rect 8668 43930 8720 43936
rect 8576 43376 8628 43382
rect 8576 43318 8628 43324
rect 8300 43104 8352 43110
rect 8300 43046 8352 43052
rect 8312 42906 8340 43046
rect 8300 42900 8352 42906
rect 8300 42842 8352 42848
rect 8588 42226 8616 43318
rect 8680 43314 8708 43930
rect 8956 43790 8984 44814
rect 8944 43784 8996 43790
rect 8944 43726 8996 43732
rect 8668 43308 8720 43314
rect 8668 43250 8720 43256
rect 8680 42294 8708 43250
rect 9036 42764 9088 42770
rect 9036 42706 9088 42712
rect 8668 42288 8720 42294
rect 8668 42230 8720 42236
rect 8392 42220 8444 42226
rect 8392 42162 8444 42168
rect 8576 42220 8628 42226
rect 8576 42162 8628 42168
rect 7932 42016 7984 42022
rect 7932 41958 7984 41964
rect 7944 41414 7972 41958
rect 7852 41386 7972 41414
rect 7748 40520 7800 40526
rect 7748 40462 7800 40468
rect 7760 40050 7788 40462
rect 7748 40044 7800 40050
rect 7748 39986 7800 39992
rect 7852 38842 7880 41386
rect 8404 41274 8432 42162
rect 8484 42152 8536 42158
rect 8484 42094 8536 42100
rect 8392 41268 8444 41274
rect 8392 41210 8444 41216
rect 8300 41200 8352 41206
rect 8496 41154 8524 42094
rect 8300 41142 8352 41148
rect 8116 41132 8168 41138
rect 8116 41074 8168 41080
rect 7932 40384 7984 40390
rect 7932 40326 7984 40332
rect 7944 40050 7972 40326
rect 8128 40186 8156 41074
rect 8312 40730 8340 41142
rect 8404 41138 8524 41154
rect 8588 41138 8616 42162
rect 8392 41132 8524 41138
rect 8444 41126 8524 41132
rect 8576 41132 8628 41138
rect 8392 41074 8444 41080
rect 8576 41074 8628 41080
rect 8404 40730 8432 41074
rect 8300 40724 8352 40730
rect 8300 40666 8352 40672
rect 8392 40724 8444 40730
rect 8392 40666 8444 40672
rect 8300 40452 8352 40458
rect 8300 40394 8352 40400
rect 8116 40180 8168 40186
rect 8116 40122 8168 40128
rect 8024 40112 8076 40118
rect 8312 40066 8340 40394
rect 8076 40060 8340 40066
rect 8024 40054 8340 40060
rect 8760 40112 8812 40118
rect 8760 40054 8812 40060
rect 7932 40044 7984 40050
rect 8036 40038 8340 40054
rect 7932 39986 7984 39992
rect 7944 39370 7972 39986
rect 8116 39840 8168 39846
rect 8116 39782 8168 39788
rect 8128 39438 8156 39782
rect 8116 39432 8168 39438
rect 8116 39374 8168 39380
rect 7932 39364 7984 39370
rect 7932 39306 7984 39312
rect 7944 39098 7972 39306
rect 7932 39092 7984 39098
rect 7932 39034 7984 39040
rect 8024 38888 8076 38894
rect 7852 38814 7972 38842
rect 8024 38830 8076 38836
rect 7840 38752 7892 38758
rect 7840 38694 7892 38700
rect 7748 37868 7800 37874
rect 7748 37810 7800 37816
rect 7484 31726 7696 31754
rect 7484 31090 7512 31726
rect 7484 31062 7696 31090
rect 7300 30790 7420 30818
rect 7300 30734 7328 30790
rect 7288 30728 7340 30734
rect 7288 30670 7340 30676
rect 6828 30660 6880 30666
rect 6828 30602 6880 30608
rect 7196 30660 7248 30666
rect 7196 30602 7248 30608
rect 6880 30492 7188 30512
rect 6880 30490 6886 30492
rect 6942 30490 6966 30492
rect 7022 30490 7046 30492
rect 7102 30490 7126 30492
rect 7182 30490 7188 30492
rect 6942 30438 6944 30490
rect 7124 30438 7126 30490
rect 6880 30436 6886 30438
rect 6942 30436 6966 30438
rect 7022 30436 7046 30438
rect 7102 30436 7126 30438
rect 7182 30436 7188 30438
rect 6880 30416 7188 30436
rect 7300 30258 7328 30670
rect 7380 30660 7432 30666
rect 7380 30602 7432 30608
rect 7288 30252 7340 30258
rect 7288 30194 7340 30200
rect 6276 29640 6328 29646
rect 6276 29582 6328 29588
rect 6288 28762 6316 29582
rect 6880 29404 7188 29424
rect 6880 29402 6886 29404
rect 6942 29402 6966 29404
rect 7022 29402 7046 29404
rect 7102 29402 7126 29404
rect 7182 29402 7188 29404
rect 6942 29350 6944 29402
rect 7124 29350 7126 29402
rect 6880 29348 6886 29350
rect 6942 29348 6966 29350
rect 7022 29348 7046 29350
rect 7102 29348 7126 29350
rect 7182 29348 7188 29350
rect 6880 29328 7188 29348
rect 6276 28756 6328 28762
rect 6276 28698 6328 28704
rect 6880 28316 7188 28336
rect 6880 28314 6886 28316
rect 6942 28314 6966 28316
rect 7022 28314 7046 28316
rect 7102 28314 7126 28316
rect 7182 28314 7188 28316
rect 6942 28262 6944 28314
rect 7124 28262 7126 28314
rect 6880 28260 6886 28262
rect 6942 28260 6966 28262
rect 7022 28260 7046 28262
rect 7102 28260 7126 28262
rect 7182 28260 7188 28262
rect 6880 28240 7188 28260
rect 7300 27402 7328 30194
rect 7392 28558 7420 30602
rect 7380 28552 7432 28558
rect 7432 28500 7512 28506
rect 7380 28494 7512 28500
rect 7392 28478 7512 28494
rect 7380 28416 7432 28422
rect 7380 28358 7432 28364
rect 7288 27396 7340 27402
rect 7288 27338 7340 27344
rect 6880 27228 7188 27248
rect 6880 27226 6886 27228
rect 6942 27226 6966 27228
rect 7022 27226 7046 27228
rect 7102 27226 7126 27228
rect 7182 27226 7188 27228
rect 6942 27174 6944 27226
rect 7124 27174 7126 27226
rect 6880 27172 6886 27174
rect 6942 27172 6966 27174
rect 7022 27172 7046 27174
rect 7102 27172 7126 27174
rect 7182 27172 7188 27174
rect 6880 27152 7188 27172
rect 7300 27062 7328 27338
rect 7392 27334 7420 28358
rect 7484 28014 7512 28478
rect 7564 28212 7616 28218
rect 7564 28154 7616 28160
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7472 27872 7524 27878
rect 7472 27814 7524 27820
rect 7380 27328 7432 27334
rect 7380 27270 7432 27276
rect 7288 27056 7340 27062
rect 7288 26998 7340 27004
rect 7300 26450 7328 26998
rect 7484 26858 7512 27814
rect 7472 26852 7524 26858
rect 7472 26794 7524 26800
rect 7484 26738 7512 26794
rect 7392 26710 7512 26738
rect 7288 26444 7340 26450
rect 7288 26386 7340 26392
rect 7392 26382 7420 26710
rect 7576 26382 7604 28154
rect 7380 26376 7432 26382
rect 7380 26318 7432 26324
rect 7564 26376 7616 26382
rect 7564 26318 7616 26324
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6380 26042 6408 26250
rect 6880 26140 7188 26160
rect 6880 26138 6886 26140
rect 6942 26138 6966 26140
rect 7022 26138 7046 26140
rect 7102 26138 7126 26140
rect 7182 26138 7188 26140
rect 6942 26086 6944 26138
rect 7124 26086 7126 26138
rect 6880 26084 6886 26086
rect 6942 26084 6966 26086
rect 7022 26084 7046 26086
rect 7102 26084 7126 26086
rect 7182 26084 7188 26086
rect 6880 26064 7188 26084
rect 6368 26036 6420 26042
rect 6368 25978 6420 25984
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 6932 25498 6960 25774
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6880 25052 7188 25072
rect 6880 25050 6886 25052
rect 6942 25050 6966 25052
rect 7022 25050 7046 25052
rect 7102 25050 7126 25052
rect 7182 25050 7188 25052
rect 6942 24998 6944 25050
rect 7124 24998 7126 25050
rect 6880 24996 6886 24998
rect 6942 24996 6966 24998
rect 7022 24996 7046 24998
rect 7102 24996 7126 24998
rect 7182 24996 7188 24998
rect 6880 24976 7188 24996
rect 6880 23964 7188 23984
rect 6880 23962 6886 23964
rect 6942 23962 6966 23964
rect 7022 23962 7046 23964
rect 7102 23962 7126 23964
rect 7182 23962 7188 23964
rect 6942 23910 6944 23962
rect 7124 23910 7126 23962
rect 6880 23908 6886 23910
rect 6942 23908 6966 23910
rect 7022 23908 7046 23910
rect 7102 23908 7126 23910
rect 7182 23908 7188 23910
rect 6880 23888 7188 23908
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 6144 23004 6224 23032
rect 6092 22986 6144 22992
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 6012 22098 6040 22918
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 6104 20482 6132 22986
rect 6368 22976 6420 22982
rect 6368 22918 6420 22924
rect 6380 22778 6408 22918
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6184 21412 6236 21418
rect 6184 21354 6236 21360
rect 6196 21010 6224 21354
rect 6472 21010 6500 23054
rect 6748 21894 6776 23598
rect 7208 23100 7236 23666
rect 7300 23662 7328 25910
rect 7392 25906 7420 26318
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 7576 25838 7604 26318
rect 7564 25832 7616 25838
rect 7564 25774 7616 25780
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 7564 23520 7616 23526
rect 7564 23462 7616 23468
rect 7288 23112 7340 23118
rect 7208 23072 7288 23100
rect 7340 23072 7420 23100
rect 7288 23054 7340 23060
rect 6880 22876 7188 22896
rect 6880 22874 6886 22876
rect 6942 22874 6966 22876
rect 7022 22874 7046 22876
rect 7102 22874 7126 22876
rect 7182 22874 7188 22876
rect 6942 22822 6944 22874
rect 7124 22822 7126 22874
rect 6880 22820 6886 22822
rect 6942 22820 6966 22822
rect 7022 22820 7046 22822
rect 7102 22820 7126 22822
rect 7182 22820 7188 22822
rect 6880 22800 7188 22820
rect 7392 22574 7420 23072
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7392 21894 7420 22510
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 6880 21788 7188 21808
rect 6880 21786 6886 21788
rect 6942 21786 6966 21788
rect 7022 21786 7046 21788
rect 7102 21786 7126 21788
rect 7182 21786 7188 21788
rect 6942 21734 6944 21786
rect 7124 21734 7126 21786
rect 6880 21732 6886 21734
rect 6942 21732 6966 21734
rect 7022 21732 7046 21734
rect 7102 21732 7126 21734
rect 7182 21732 7188 21734
rect 6880 21712 7188 21732
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6012 20454 6132 20482
rect 6472 20466 6500 20946
rect 7392 20942 7420 21830
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 6880 20700 7188 20720
rect 6880 20698 6886 20700
rect 6942 20698 6966 20700
rect 7022 20698 7046 20700
rect 7102 20698 7126 20700
rect 7182 20698 7188 20700
rect 6942 20646 6944 20698
rect 7124 20646 7126 20698
rect 6880 20644 6886 20646
rect 6942 20644 6966 20646
rect 7022 20644 7046 20646
rect 7102 20644 7126 20646
rect 7182 20644 7188 20646
rect 6880 20624 7188 20644
rect 7392 20466 7420 20878
rect 7484 20602 7512 21490
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 6460 20460 6512 20466
rect 6012 20262 6040 20454
rect 6460 20402 6512 20408
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5908 17808 5960 17814
rect 5908 17750 5960 17756
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16114 5764 16390
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5276 15094 5304 15642
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4448 14346 4476 14962
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 3915 13628 4223 13648
rect 3915 13626 3921 13628
rect 3977 13626 4001 13628
rect 4057 13626 4081 13628
rect 4137 13626 4161 13628
rect 4217 13626 4223 13628
rect 3977 13574 3979 13626
rect 4159 13574 4161 13626
rect 3915 13572 3921 13574
rect 3977 13572 4001 13574
rect 4057 13572 4081 13574
rect 4137 13572 4161 13574
rect 4217 13572 4223 13574
rect 3915 13552 4223 13572
rect 3915 12540 4223 12560
rect 3915 12538 3921 12540
rect 3977 12538 4001 12540
rect 4057 12538 4081 12540
rect 4137 12538 4161 12540
rect 4217 12538 4223 12540
rect 3977 12486 3979 12538
rect 4159 12486 4161 12538
rect 3915 12484 3921 12486
rect 3977 12484 4001 12486
rect 4057 12484 4081 12486
rect 4137 12484 4161 12486
rect 4217 12484 4223 12486
rect 3915 12464 4223 12484
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3804 11150 3832 12174
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 3915 11452 4223 11472
rect 3915 11450 3921 11452
rect 3977 11450 4001 11452
rect 4057 11450 4081 11452
rect 4137 11450 4161 11452
rect 4217 11450 4223 11452
rect 3977 11398 3979 11450
rect 4159 11398 4161 11450
rect 3915 11396 3921 11398
rect 3977 11396 4001 11398
rect 4057 11396 4081 11398
rect 4137 11396 4161 11398
rect 4217 11396 4223 11398
rect 3915 11376 4223 11396
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 1400 8968 1452 8974
rect 1398 8936 1400 8945
rect 1452 8936 1454 8945
rect 1398 8871 1454 8880
rect 3804 8498 3832 11086
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4264 10742 4292 11018
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4448 10674 4476 11494
rect 5000 11286 5028 11698
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 3915 10364 4223 10384
rect 3915 10362 3921 10364
rect 3977 10362 4001 10364
rect 4057 10362 4081 10364
rect 4137 10362 4161 10364
rect 4217 10362 4223 10364
rect 3977 10310 3979 10362
rect 4159 10310 4161 10362
rect 3915 10308 3921 10310
rect 3977 10308 4001 10310
rect 4057 10308 4081 10310
rect 4137 10308 4161 10310
rect 4217 10308 4223 10310
rect 3915 10288 4223 10308
rect 3915 9276 4223 9296
rect 3915 9274 3921 9276
rect 3977 9274 4001 9276
rect 4057 9274 4081 9276
rect 4137 9274 4161 9276
rect 4217 9274 4223 9276
rect 3977 9222 3979 9274
rect 4159 9222 4161 9274
rect 3915 9220 3921 9222
rect 3977 9220 4001 9222
rect 4057 9220 4081 9222
rect 4137 9220 4161 9222
rect 4217 9220 4223 9222
rect 3915 9200 4223 9220
rect 4632 9042 4660 10474
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 9178 4752 9318
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4816 8974 4844 10610
rect 5000 9586 5028 11222
rect 5092 11082 5120 11698
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5092 10062 5120 11018
rect 5552 10130 5580 11698
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 10606 5672 11494
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5828 10674 5856 10950
rect 5920 10674 5948 11698
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5828 10198 5856 10610
rect 5920 10266 5948 10610
rect 6012 10538 6040 20198
rect 6880 19612 7188 19632
rect 6880 19610 6886 19612
rect 6942 19610 6966 19612
rect 7022 19610 7046 19612
rect 7102 19610 7126 19612
rect 7182 19610 7188 19612
rect 6942 19558 6944 19610
rect 7124 19558 7126 19610
rect 6880 19556 6886 19558
rect 6942 19556 6966 19558
rect 7022 19556 7046 19558
rect 7102 19556 7126 19558
rect 7182 19556 7188 19558
rect 6880 19536 7188 19556
rect 6880 18524 7188 18544
rect 6880 18522 6886 18524
rect 6942 18522 6966 18524
rect 7022 18522 7046 18524
rect 7102 18522 7126 18524
rect 7182 18522 7188 18524
rect 6942 18470 6944 18522
rect 7124 18470 7126 18522
rect 6880 18468 6886 18470
rect 6942 18468 6966 18470
rect 7022 18468 7046 18470
rect 7102 18468 7126 18470
rect 7182 18468 7188 18470
rect 6880 18448 7188 18468
rect 6368 18352 6420 18358
rect 6368 18294 6420 18300
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6196 16182 6224 17682
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6288 16726 6316 17614
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6104 15473 6132 15914
rect 6196 15502 6224 16118
rect 6184 15496 6236 15502
rect 6090 15464 6146 15473
rect 6184 15438 6236 15444
rect 6090 15399 6092 15408
rect 6144 15399 6146 15408
rect 6092 15370 6144 15376
rect 6288 11626 6316 16662
rect 6380 16590 6408 18294
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6472 15706 6500 17614
rect 6564 15910 6592 18226
rect 6748 17746 6776 18226
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 6920 18080 6972 18086
rect 6840 18028 6920 18034
rect 6840 18022 6972 18028
rect 6840 18006 6960 18022
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6644 17536 6696 17542
rect 6840 17524 6868 18006
rect 7208 17882 7236 18090
rect 7196 17876 7248 17882
rect 7576 17864 7604 23462
rect 7668 22642 7696 31062
rect 7760 30666 7788 37810
rect 7852 37194 7880 38694
rect 7944 37398 7972 38814
rect 8036 37806 8064 38830
rect 8128 38418 8156 39374
rect 8208 38956 8260 38962
rect 8208 38898 8260 38904
rect 8116 38412 8168 38418
rect 8116 38354 8168 38360
rect 8220 38010 8248 38898
rect 8208 38004 8260 38010
rect 8208 37946 8260 37952
rect 8312 37806 8340 40038
rect 8484 39296 8536 39302
rect 8484 39238 8536 39244
rect 8496 38978 8524 39238
rect 8404 38962 8524 38978
rect 8772 38962 8800 40054
rect 8944 40044 8996 40050
rect 8944 39986 8996 39992
rect 8956 39098 8984 39986
rect 8944 39092 8996 39098
rect 8944 39034 8996 39040
rect 8392 38956 8524 38962
rect 8444 38950 8524 38956
rect 8760 38956 8812 38962
rect 8392 38898 8444 38904
rect 8760 38898 8812 38904
rect 8772 37942 8800 38898
rect 8760 37936 8812 37942
rect 8760 37878 8812 37884
rect 8852 37868 8904 37874
rect 8852 37810 8904 37816
rect 8024 37800 8076 37806
rect 8024 37742 8076 37748
rect 8300 37800 8352 37806
rect 8300 37742 8352 37748
rect 7932 37392 7984 37398
rect 7932 37334 7984 37340
rect 7840 37188 7892 37194
rect 7840 37130 7892 37136
rect 7932 37120 7984 37126
rect 7932 37062 7984 37068
rect 7840 36780 7892 36786
rect 7840 36722 7892 36728
rect 7852 36378 7880 36722
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 7944 36174 7972 37062
rect 7932 36168 7984 36174
rect 7932 36110 7984 36116
rect 8036 34202 8064 37742
rect 8208 37392 8260 37398
rect 8208 37334 8260 37340
rect 8116 36848 8168 36854
rect 8116 36790 8168 36796
rect 8128 36242 8156 36790
rect 8116 36236 8168 36242
rect 8116 36178 8168 36184
rect 8024 34196 8076 34202
rect 8024 34138 8076 34144
rect 8220 34082 8248 37334
rect 8300 37188 8352 37194
rect 8300 37130 8352 37136
rect 8312 36174 8340 37130
rect 8392 36304 8444 36310
rect 8392 36246 8444 36252
rect 8300 36168 8352 36174
rect 8300 36110 8352 36116
rect 7944 34054 8248 34082
rect 7944 33153 7972 34054
rect 8024 33924 8076 33930
rect 8024 33866 8076 33872
rect 7930 33144 7986 33153
rect 7930 33079 7986 33088
rect 7932 32496 7984 32502
rect 7932 32438 7984 32444
rect 7944 31822 7972 32438
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 7840 31680 7892 31686
rect 7840 31622 7892 31628
rect 7852 31278 7880 31622
rect 7840 31272 7892 31278
rect 7840 31214 7892 31220
rect 7748 30660 7800 30666
rect 7748 30602 7800 30608
rect 7852 30598 7880 31214
rect 7944 31142 7972 31758
rect 8036 31754 8064 33866
rect 8312 33590 8340 36110
rect 8404 35630 8432 36246
rect 8864 36038 8892 37810
rect 8852 36032 8904 36038
rect 8852 35974 8904 35980
rect 8864 35698 8892 35974
rect 8852 35692 8904 35698
rect 8852 35634 8904 35640
rect 8392 35624 8444 35630
rect 8392 35566 8444 35572
rect 8300 33584 8352 33590
rect 8300 33526 8352 33532
rect 8116 33516 8168 33522
rect 8116 33458 8168 33464
rect 8208 33516 8260 33522
rect 8208 33458 8260 33464
rect 8128 32842 8156 33458
rect 8220 33130 8248 33458
rect 8312 33266 8340 33526
rect 8760 33380 8812 33386
rect 8760 33322 8812 33328
rect 8312 33238 8432 33266
rect 8220 33114 8340 33130
rect 8220 33108 8352 33114
rect 8220 33102 8300 33108
rect 8300 33050 8352 33056
rect 8208 32972 8260 32978
rect 8208 32914 8260 32920
rect 8116 32836 8168 32842
rect 8116 32778 8168 32784
rect 8128 32434 8156 32778
rect 8116 32428 8168 32434
rect 8116 32370 8168 32376
rect 8220 32366 8248 32914
rect 8208 32360 8260 32366
rect 8312 32348 8340 33050
rect 8404 32910 8432 33238
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 8404 32502 8432 32846
rect 8392 32496 8444 32502
rect 8392 32438 8444 32444
rect 8392 32360 8444 32366
rect 8312 32320 8392 32348
rect 8208 32302 8260 32308
rect 8392 32302 8444 32308
rect 8036 31726 8156 31754
rect 7932 31136 7984 31142
rect 7932 31078 7984 31084
rect 7840 30592 7892 30598
rect 7840 30534 7892 30540
rect 7852 29714 7880 30534
rect 7840 29708 7892 29714
rect 7840 29650 7892 29656
rect 7840 28552 7892 28558
rect 7840 28494 7892 28500
rect 7852 28218 7880 28494
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 8024 27872 8076 27878
rect 8024 27814 8076 27820
rect 8036 26586 8064 27814
rect 8024 26580 8076 26586
rect 8024 26522 8076 26528
rect 8036 26382 8064 26522
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 8128 23594 8156 31726
rect 8220 28014 8248 32302
rect 8300 31136 8352 31142
rect 8300 31078 8352 31084
rect 8312 30326 8340 31078
rect 8404 30938 8432 32302
rect 8772 31346 8800 33322
rect 8944 33312 8996 33318
rect 8944 33254 8996 33260
rect 8956 33114 8984 33254
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 9048 32978 9076 42706
rect 9140 42566 9168 45902
rect 9220 45824 9272 45830
rect 9220 45766 9272 45772
rect 9232 43790 9260 45766
rect 12811 45724 13119 45744
rect 12811 45722 12817 45724
rect 12873 45722 12897 45724
rect 12953 45722 12977 45724
rect 13033 45722 13057 45724
rect 13113 45722 13119 45724
rect 12873 45670 12875 45722
rect 13055 45670 13057 45722
rect 12811 45668 12817 45670
rect 12873 45668 12897 45670
rect 12953 45668 12977 45670
rect 13033 45668 13057 45670
rect 13113 45668 13119 45670
rect 12811 45648 13119 45668
rect 10324 45552 10376 45558
rect 10324 45494 10376 45500
rect 10232 45280 10284 45286
rect 10232 45222 10284 45228
rect 9846 45180 10154 45200
rect 9846 45178 9852 45180
rect 9908 45178 9932 45180
rect 9988 45178 10012 45180
rect 10068 45178 10092 45180
rect 10148 45178 10154 45180
rect 9908 45126 9910 45178
rect 10090 45126 10092 45178
rect 9846 45124 9852 45126
rect 9908 45124 9932 45126
rect 9988 45124 10012 45126
rect 10068 45124 10092 45126
rect 10148 45124 10154 45126
rect 9846 45104 10154 45124
rect 9772 44192 9824 44198
rect 9772 44134 9824 44140
rect 9220 43784 9272 43790
rect 9220 43726 9272 43732
rect 9220 43308 9272 43314
rect 9220 43250 9272 43256
rect 9680 43308 9732 43314
rect 9680 43250 9732 43256
rect 9128 42560 9180 42566
rect 9128 42502 9180 42508
rect 9232 42362 9260 43250
rect 9588 43172 9640 43178
rect 9588 43114 9640 43120
rect 9600 42566 9628 43114
rect 9692 42702 9720 43250
rect 9784 42702 9812 44134
rect 9846 44092 10154 44112
rect 9846 44090 9852 44092
rect 9908 44090 9932 44092
rect 9988 44090 10012 44092
rect 10068 44090 10092 44092
rect 10148 44090 10154 44092
rect 9908 44038 9910 44090
rect 10090 44038 10092 44090
rect 9846 44036 9852 44038
rect 9908 44036 9932 44038
rect 9988 44036 10012 44038
rect 10068 44036 10092 44038
rect 10148 44036 10154 44038
rect 9846 44016 10154 44036
rect 10244 43994 10272 45222
rect 10336 44742 10364 45494
rect 10416 45484 10468 45490
rect 10416 45426 10468 45432
rect 11520 45484 11572 45490
rect 11520 45426 11572 45432
rect 12072 45484 12124 45490
rect 12072 45426 12124 45432
rect 10428 44810 10456 45426
rect 10876 44872 10928 44878
rect 10876 44814 10928 44820
rect 11428 44872 11480 44878
rect 11428 44814 11480 44820
rect 10416 44804 10468 44810
rect 10416 44746 10468 44752
rect 10888 44742 10916 44814
rect 11336 44804 11388 44810
rect 11336 44746 11388 44752
rect 10324 44736 10376 44742
rect 10324 44678 10376 44684
rect 10876 44736 10928 44742
rect 10876 44678 10928 44684
rect 10324 44396 10376 44402
rect 10324 44338 10376 44344
rect 10232 43988 10284 43994
rect 10232 43930 10284 43936
rect 10244 43722 10272 43930
rect 10232 43716 10284 43722
rect 10232 43658 10284 43664
rect 10244 43246 10272 43658
rect 10336 43382 10364 44338
rect 10888 43858 10916 44678
rect 10876 43852 10928 43858
rect 10876 43794 10928 43800
rect 11348 43790 11376 44746
rect 11440 43994 11468 44814
rect 11428 43988 11480 43994
rect 11428 43930 11480 43936
rect 10784 43784 10836 43790
rect 10784 43726 10836 43732
rect 11336 43784 11388 43790
rect 11336 43726 11388 43732
rect 10796 43450 10824 43726
rect 10968 43648 11020 43654
rect 10968 43590 11020 43596
rect 10784 43444 10836 43450
rect 10784 43386 10836 43392
rect 10980 43382 11008 43590
rect 10324 43376 10376 43382
rect 10324 43318 10376 43324
rect 10968 43376 11020 43382
rect 10968 43318 11020 43324
rect 10784 43308 10836 43314
rect 10784 43250 10836 43256
rect 10232 43240 10284 43246
rect 10232 43182 10284 43188
rect 10508 43104 10560 43110
rect 10508 43046 10560 43052
rect 9846 43004 10154 43024
rect 9846 43002 9852 43004
rect 9908 43002 9932 43004
rect 9988 43002 10012 43004
rect 10068 43002 10092 43004
rect 10148 43002 10154 43004
rect 9908 42950 9910 43002
rect 10090 42950 10092 43002
rect 9846 42948 9852 42950
rect 9908 42948 9932 42950
rect 9988 42948 10012 42950
rect 10068 42948 10092 42950
rect 10148 42948 10154 42950
rect 9846 42928 10154 42948
rect 9680 42696 9732 42702
rect 9680 42638 9732 42644
rect 9772 42696 9824 42702
rect 9772 42638 9824 42644
rect 9588 42560 9640 42566
rect 9588 42502 9640 42508
rect 9220 42356 9272 42362
rect 9220 42298 9272 42304
rect 9600 42226 9628 42502
rect 9784 42226 9812 42638
rect 10520 42362 10548 43046
rect 10508 42356 10560 42362
rect 10508 42298 10560 42304
rect 9588 42220 9640 42226
rect 9588 42162 9640 42168
rect 9772 42220 9824 42226
rect 9772 42162 9824 42168
rect 9680 40520 9732 40526
rect 9680 40462 9732 40468
rect 9692 39642 9720 40462
rect 9680 39636 9732 39642
rect 9680 39578 9732 39584
rect 9692 38962 9720 39578
rect 9784 39370 9812 42162
rect 9846 41916 10154 41936
rect 9846 41914 9852 41916
rect 9908 41914 9932 41916
rect 9988 41914 10012 41916
rect 10068 41914 10092 41916
rect 10148 41914 10154 41916
rect 9908 41862 9910 41914
rect 10090 41862 10092 41914
rect 9846 41860 9852 41862
rect 9908 41860 9932 41862
rect 9988 41860 10012 41862
rect 10068 41860 10092 41862
rect 10148 41860 10154 41862
rect 9846 41840 10154 41860
rect 9846 40828 10154 40848
rect 9846 40826 9852 40828
rect 9908 40826 9932 40828
rect 9988 40826 10012 40828
rect 10068 40826 10092 40828
rect 10148 40826 10154 40828
rect 9908 40774 9910 40826
rect 10090 40774 10092 40826
rect 9846 40772 9852 40774
rect 9908 40772 9932 40774
rect 9988 40772 10012 40774
rect 10068 40772 10092 40774
rect 10148 40772 10154 40774
rect 9846 40752 10154 40772
rect 10232 40044 10284 40050
rect 10232 39986 10284 39992
rect 9846 39740 10154 39760
rect 9846 39738 9852 39740
rect 9908 39738 9932 39740
rect 9988 39738 10012 39740
rect 10068 39738 10092 39740
rect 10148 39738 10154 39740
rect 9908 39686 9910 39738
rect 10090 39686 10092 39738
rect 9846 39684 9852 39686
rect 9908 39684 9932 39686
rect 9988 39684 10012 39686
rect 10068 39684 10092 39686
rect 10148 39684 10154 39686
rect 9846 39664 10154 39684
rect 10244 39574 10272 39986
rect 10324 39976 10376 39982
rect 10324 39918 10376 39924
rect 10232 39568 10284 39574
rect 10232 39510 10284 39516
rect 9956 39500 10008 39506
rect 9876 39460 9956 39488
rect 9772 39364 9824 39370
rect 9772 39306 9824 39312
rect 9680 38956 9732 38962
rect 9680 38898 9732 38904
rect 9692 38350 9720 38898
rect 9876 38842 9904 39460
rect 9956 39442 10008 39448
rect 10244 38894 10272 39510
rect 9784 38814 9904 38842
rect 10232 38888 10284 38894
rect 10232 38830 10284 38836
rect 10336 38826 10364 39918
rect 10796 39846 10824 43250
rect 10876 43104 10928 43110
rect 10876 43046 10928 43052
rect 10888 42650 10916 43046
rect 10980 42770 11008 43318
rect 10968 42764 11020 42770
rect 10968 42706 11020 42712
rect 10888 42622 11008 42650
rect 10876 42220 10928 42226
rect 10876 42162 10928 42168
rect 10784 39840 10836 39846
rect 10784 39782 10836 39788
rect 10888 39386 10916 42162
rect 10704 39358 10916 39386
rect 10416 39296 10468 39302
rect 10416 39238 10468 39244
rect 10428 38962 10456 39238
rect 10508 39024 10560 39030
rect 10508 38966 10560 38972
rect 10416 38956 10468 38962
rect 10416 38898 10468 38904
rect 10324 38820 10376 38826
rect 9784 38418 9812 38814
rect 10324 38762 10376 38768
rect 9846 38652 10154 38672
rect 9846 38650 9852 38652
rect 9908 38650 9932 38652
rect 9988 38650 10012 38652
rect 10068 38650 10092 38652
rect 10148 38650 10154 38652
rect 9908 38598 9910 38650
rect 10090 38598 10092 38650
rect 9846 38596 9852 38598
rect 9908 38596 9932 38598
rect 9988 38596 10012 38598
rect 10068 38596 10092 38598
rect 10148 38596 10154 38598
rect 9846 38576 10154 38596
rect 9772 38412 9824 38418
rect 9772 38354 9824 38360
rect 10324 38412 10376 38418
rect 10324 38354 10376 38360
rect 9680 38344 9732 38350
rect 9680 38286 9732 38292
rect 10232 38344 10284 38350
rect 10232 38286 10284 38292
rect 9680 38004 9732 38010
rect 9680 37946 9732 37952
rect 9404 37664 9456 37670
rect 9404 37606 9456 37612
rect 9128 37256 9180 37262
rect 9128 37198 9180 37204
rect 9140 34082 9168 37198
rect 9416 36786 9444 37606
rect 9404 36780 9456 36786
rect 9404 36722 9456 36728
rect 9220 36100 9272 36106
rect 9220 36042 9272 36048
rect 9232 35834 9260 36042
rect 9220 35828 9272 35834
rect 9220 35770 9272 35776
rect 9404 35692 9456 35698
rect 9404 35634 9456 35640
rect 9588 35692 9640 35698
rect 9588 35634 9640 35640
rect 9140 34054 9260 34082
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 9036 32972 9088 32978
rect 9036 32914 9088 32920
rect 9140 32910 9168 33934
rect 9232 33454 9260 34054
rect 9220 33448 9272 33454
rect 9220 33390 9272 33396
rect 9128 32904 9180 32910
rect 9128 32846 9180 32852
rect 8852 32564 8904 32570
rect 8852 32506 8904 32512
rect 8760 31340 8812 31346
rect 8760 31282 8812 31288
rect 8864 31278 8892 32506
rect 9140 31414 9168 32846
rect 9416 31890 9444 35634
rect 9600 32026 9628 35634
rect 9692 35630 9720 37946
rect 9772 37868 9824 37874
rect 9772 37810 9824 37816
rect 9784 37398 9812 37810
rect 10244 37806 10272 38286
rect 10232 37800 10284 37806
rect 10232 37742 10284 37748
rect 9846 37564 10154 37584
rect 9846 37562 9852 37564
rect 9908 37562 9932 37564
rect 9988 37562 10012 37564
rect 10068 37562 10092 37564
rect 10148 37562 10154 37564
rect 9908 37510 9910 37562
rect 10090 37510 10092 37562
rect 9846 37508 9852 37510
rect 9908 37508 9932 37510
rect 9988 37508 10012 37510
rect 10068 37508 10092 37510
rect 10148 37508 10154 37510
rect 9846 37488 10154 37508
rect 9772 37392 9824 37398
rect 9772 37334 9824 37340
rect 10244 36922 10272 37742
rect 10232 36916 10284 36922
rect 10232 36858 10284 36864
rect 9846 36476 10154 36496
rect 9846 36474 9852 36476
rect 9908 36474 9932 36476
rect 9988 36474 10012 36476
rect 10068 36474 10092 36476
rect 10148 36474 10154 36476
rect 9908 36422 9910 36474
rect 10090 36422 10092 36474
rect 9846 36420 9852 36422
rect 9908 36420 9932 36422
rect 9988 36420 10012 36422
rect 10068 36420 10092 36422
rect 10148 36420 10154 36422
rect 9846 36400 10154 36420
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 9692 33046 9720 35566
rect 9846 35388 10154 35408
rect 9846 35386 9852 35388
rect 9908 35386 9932 35388
rect 9988 35386 10012 35388
rect 10068 35386 10092 35388
rect 10148 35386 10154 35388
rect 9908 35334 9910 35386
rect 10090 35334 10092 35386
rect 9846 35332 9852 35334
rect 9908 35332 9932 35334
rect 9988 35332 10012 35334
rect 10068 35332 10092 35334
rect 10148 35332 10154 35334
rect 9846 35312 10154 35332
rect 9846 34300 10154 34320
rect 9846 34298 9852 34300
rect 9908 34298 9932 34300
rect 9988 34298 10012 34300
rect 10068 34298 10092 34300
rect 10148 34298 10154 34300
rect 9908 34246 9910 34298
rect 10090 34246 10092 34298
rect 9846 34244 9852 34246
rect 9908 34244 9932 34246
rect 9988 34244 10012 34246
rect 10068 34244 10092 34246
rect 10148 34244 10154 34246
rect 9846 34224 10154 34244
rect 10232 33312 10284 33318
rect 10232 33254 10284 33260
rect 9846 33212 10154 33232
rect 9846 33210 9852 33212
rect 9908 33210 9932 33212
rect 9988 33210 10012 33212
rect 10068 33210 10092 33212
rect 10148 33210 10154 33212
rect 9908 33158 9910 33210
rect 10090 33158 10092 33210
rect 9846 33156 9852 33158
rect 9908 33156 9932 33158
rect 9988 33156 10012 33158
rect 10068 33156 10092 33158
rect 10148 33156 10154 33158
rect 9846 33136 10154 33156
rect 9680 33040 9732 33046
rect 9732 33000 9812 33028
rect 9680 32982 9732 32988
rect 9680 32496 9732 32502
rect 9680 32438 9732 32444
rect 9588 32020 9640 32026
rect 9588 31962 9640 31968
rect 9404 31884 9456 31890
rect 9404 31826 9456 31832
rect 9128 31408 9180 31414
rect 9128 31350 9180 31356
rect 8852 31272 8904 31278
rect 8852 31214 8904 31220
rect 8392 30932 8444 30938
rect 8392 30874 8444 30880
rect 9140 30818 9168 31350
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 9048 30790 9168 30818
rect 9048 30734 9076 30790
rect 9600 30734 9628 31214
rect 9036 30728 9088 30734
rect 9036 30670 9088 30676
rect 9588 30728 9640 30734
rect 9588 30670 9640 30676
rect 9048 30394 9076 30670
rect 9036 30388 9088 30394
rect 9036 30330 9088 30336
rect 8300 30320 8352 30326
rect 8300 30262 8352 30268
rect 9600 29646 9628 30670
rect 9692 30666 9720 32438
rect 9784 31210 9812 33000
rect 10244 32978 10272 33254
rect 10232 32972 10284 32978
rect 10232 32914 10284 32920
rect 10244 32502 10272 32914
rect 10336 32570 10364 38354
rect 10416 37664 10468 37670
rect 10416 37606 10468 37612
rect 10428 37466 10456 37606
rect 10416 37460 10468 37466
rect 10416 37402 10468 37408
rect 10520 37262 10548 38966
rect 10600 38820 10652 38826
rect 10600 38762 10652 38768
rect 10612 38214 10640 38762
rect 10600 38208 10652 38214
rect 10600 38150 10652 38156
rect 10612 37874 10640 38150
rect 10704 37942 10732 39358
rect 10980 39012 11008 42622
rect 11532 42226 11560 45426
rect 12084 44878 12112 45426
rect 13268 45280 13320 45286
rect 13268 45222 13320 45228
rect 11612 44872 11664 44878
rect 11612 44814 11664 44820
rect 12072 44872 12124 44878
rect 12072 44814 12124 44820
rect 11624 43926 11652 44814
rect 12084 44538 12112 44814
rect 12811 44636 13119 44656
rect 12811 44634 12817 44636
rect 12873 44634 12897 44636
rect 12953 44634 12977 44636
rect 13033 44634 13057 44636
rect 13113 44634 13119 44636
rect 12873 44582 12875 44634
rect 13055 44582 13057 44634
rect 12811 44580 12817 44582
rect 12873 44580 12897 44582
rect 12953 44580 12977 44582
rect 13033 44580 13057 44582
rect 13113 44580 13119 44582
rect 12811 44560 13119 44580
rect 12072 44532 12124 44538
rect 12072 44474 12124 44480
rect 12808 44396 12860 44402
rect 12808 44338 12860 44344
rect 12820 43994 12848 44338
rect 12808 43988 12860 43994
rect 12808 43930 12860 43936
rect 13280 43926 13308 45222
rect 15776 45180 16084 45200
rect 15776 45178 15782 45180
rect 15838 45178 15862 45180
rect 15918 45178 15942 45180
rect 15998 45178 16022 45180
rect 16078 45178 16084 45180
rect 15838 45126 15840 45178
rect 16020 45126 16022 45178
rect 15776 45124 15782 45126
rect 15838 45124 15862 45126
rect 15918 45124 15942 45126
rect 15998 45124 16022 45126
rect 16078 45124 16084 45126
rect 15776 45104 16084 45124
rect 17880 45014 17908 46990
rect 17868 45008 17920 45014
rect 17868 44950 17920 44956
rect 13820 44396 13872 44402
rect 13820 44338 13872 44344
rect 11612 43920 11664 43926
rect 11612 43862 11664 43868
rect 13268 43920 13320 43926
rect 13268 43862 13320 43868
rect 11624 43110 11652 43862
rect 12256 43852 12308 43858
rect 12256 43794 12308 43800
rect 11980 43648 12032 43654
rect 11980 43590 12032 43596
rect 11888 43308 11940 43314
rect 11888 43250 11940 43256
rect 11612 43104 11664 43110
rect 11612 43046 11664 43052
rect 11520 42220 11572 42226
rect 11520 42162 11572 42168
rect 11704 39840 11756 39846
rect 11704 39782 11756 39788
rect 11060 39568 11112 39574
rect 11060 39510 11112 39516
rect 11072 39098 11100 39510
rect 11716 39438 11744 39782
rect 11900 39642 11928 43250
rect 11992 43246 12020 43590
rect 11980 43240 12032 43246
rect 11980 43182 12032 43188
rect 12072 40044 12124 40050
rect 12072 39986 12124 39992
rect 11888 39636 11940 39642
rect 11888 39578 11940 39584
rect 11704 39432 11756 39438
rect 11704 39374 11756 39380
rect 11796 39432 11848 39438
rect 11796 39374 11848 39380
rect 11060 39092 11112 39098
rect 11060 39034 11112 39040
rect 10796 38984 11008 39012
rect 10692 37936 10744 37942
rect 10692 37878 10744 37884
rect 10600 37868 10652 37874
rect 10600 37810 10652 37816
rect 10508 37256 10560 37262
rect 10508 37198 10560 37204
rect 10520 36378 10548 37198
rect 10508 36372 10560 36378
rect 10508 36314 10560 36320
rect 10612 36174 10640 37810
rect 10692 37800 10744 37806
rect 10692 37742 10744 37748
rect 10704 37330 10732 37742
rect 10692 37324 10744 37330
rect 10692 37266 10744 37272
rect 10600 36168 10652 36174
rect 10600 36110 10652 36116
rect 10600 35692 10652 35698
rect 10600 35634 10652 35640
rect 10416 35012 10468 35018
rect 10416 34954 10468 34960
rect 10428 34746 10456 34954
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10508 34604 10560 34610
rect 10508 34546 10560 34552
rect 10416 33448 10468 33454
rect 10416 33390 10468 33396
rect 10428 33046 10456 33390
rect 10416 33040 10468 33046
rect 10416 32982 10468 32988
rect 10324 32564 10376 32570
rect 10324 32506 10376 32512
rect 10232 32496 10284 32502
rect 10232 32438 10284 32444
rect 9846 32124 10154 32144
rect 9846 32122 9852 32124
rect 9908 32122 9932 32124
rect 9988 32122 10012 32124
rect 10068 32122 10092 32124
rect 10148 32122 10154 32124
rect 9908 32070 9910 32122
rect 10090 32070 10092 32122
rect 9846 32068 9852 32070
rect 9908 32068 9932 32070
rect 9988 32068 10012 32070
rect 10068 32068 10092 32070
rect 10148 32068 10154 32070
rect 9846 32048 10154 32068
rect 10336 31890 10364 32506
rect 10324 31884 10376 31890
rect 10324 31826 10376 31832
rect 10416 31884 10468 31890
rect 10416 31826 10468 31832
rect 10336 31754 10364 31826
rect 10428 31754 10456 31826
rect 10244 31726 10364 31754
rect 10416 31748 10468 31754
rect 9956 31680 10008 31686
rect 9956 31622 10008 31628
rect 9968 31346 9996 31622
rect 10140 31476 10192 31482
rect 10140 31418 10192 31424
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9680 30660 9732 30666
rect 9680 30602 9732 30608
rect 9692 30258 9720 30602
rect 9680 30252 9732 30258
rect 9680 30194 9732 30200
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9692 29714 9720 29990
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 8312 27674 8340 28018
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 9692 27470 9720 29514
rect 9784 27606 9812 31146
rect 10152 31124 10180 31418
rect 10244 31278 10272 31726
rect 10416 31690 10468 31696
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10232 31272 10284 31278
rect 10232 31214 10284 31220
rect 10336 31124 10364 31282
rect 10152 31096 10364 31124
rect 9846 31036 10154 31056
rect 9846 31034 9852 31036
rect 9908 31034 9932 31036
rect 9988 31034 10012 31036
rect 10068 31034 10092 31036
rect 10148 31034 10154 31036
rect 9908 30982 9910 31034
rect 10090 30982 10092 31034
rect 9846 30980 9852 30982
rect 9908 30980 9932 30982
rect 9988 30980 10012 30982
rect 10068 30980 10092 30982
rect 10148 30980 10154 30982
rect 9846 30960 10154 30980
rect 9956 30592 10008 30598
rect 9956 30534 10008 30540
rect 9968 30326 9996 30534
rect 9956 30320 10008 30326
rect 9956 30262 10008 30268
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 9846 29948 10154 29968
rect 9846 29946 9852 29948
rect 9908 29946 9932 29948
rect 9988 29946 10012 29948
rect 10068 29946 10092 29948
rect 10148 29946 10154 29948
rect 9908 29894 9910 29946
rect 10090 29894 10092 29946
rect 9846 29892 9852 29894
rect 9908 29892 9932 29894
rect 9988 29892 10012 29894
rect 10068 29892 10092 29894
rect 10148 29892 10154 29894
rect 9846 29872 10154 29892
rect 10244 29646 10272 30194
rect 10232 29640 10284 29646
rect 10232 29582 10284 29588
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 9846 28860 10154 28880
rect 9846 28858 9852 28860
rect 9908 28858 9932 28860
rect 9988 28858 10012 28860
rect 10068 28858 10092 28860
rect 10148 28858 10154 28860
rect 9908 28806 9910 28858
rect 10090 28806 10092 28858
rect 9846 28804 9852 28806
rect 9908 28804 9932 28806
rect 9988 28804 10012 28806
rect 10068 28804 10092 28806
rect 10148 28804 10154 28806
rect 9846 28784 10154 28804
rect 10244 28558 10272 29446
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 9846 27772 10154 27792
rect 9846 27770 9852 27772
rect 9908 27770 9932 27772
rect 9988 27770 10012 27772
rect 10068 27770 10092 27772
rect 10148 27770 10154 27772
rect 9908 27718 9910 27770
rect 10090 27718 10092 27770
rect 9846 27716 9852 27718
rect 9908 27716 9932 27718
rect 9988 27716 10012 27718
rect 10068 27716 10092 27718
rect 10148 27716 10154 27718
rect 9846 27696 10154 27716
rect 9772 27600 9824 27606
rect 9772 27542 9824 27548
rect 10244 27538 10272 28358
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 10336 27470 10364 31096
rect 10428 30938 10456 31690
rect 10416 30932 10468 30938
rect 10416 30874 10468 30880
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10428 30258 10456 30534
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10416 28008 10468 28014
rect 10416 27950 10468 27956
rect 10428 27606 10456 27950
rect 10416 27600 10468 27606
rect 10416 27542 10468 27548
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 10324 27464 10376 27470
rect 10324 27406 10376 27412
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9416 27062 9444 27270
rect 9692 27130 9720 27406
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9404 27056 9456 27062
rect 9404 26998 9456 27004
rect 8392 26988 8444 26994
rect 8392 26930 8444 26936
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 8404 26586 8432 26930
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 9784 26450 9812 26930
rect 9846 26684 10154 26704
rect 9846 26682 9852 26684
rect 9908 26682 9932 26684
rect 9988 26682 10012 26684
rect 10068 26682 10092 26684
rect 10148 26682 10154 26684
rect 9908 26630 9910 26682
rect 10090 26630 10092 26682
rect 9846 26628 9852 26630
rect 9908 26628 9932 26630
rect 9988 26628 10012 26630
rect 10068 26628 10092 26630
rect 10148 26628 10154 26630
rect 9846 26608 10154 26628
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8404 26042 8432 26318
rect 10336 26042 10364 27406
rect 10416 26308 10468 26314
rect 10416 26250 10468 26256
rect 10428 26042 10456 26250
rect 8392 26036 8444 26042
rect 8392 25978 8444 25984
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 9846 25596 10154 25616
rect 9846 25594 9852 25596
rect 9908 25594 9932 25596
rect 9988 25594 10012 25596
rect 10068 25594 10092 25596
rect 10148 25594 10154 25596
rect 9908 25542 9910 25594
rect 10090 25542 10092 25594
rect 9846 25540 9852 25542
rect 9908 25540 9932 25542
rect 9988 25540 10012 25542
rect 10068 25540 10092 25542
rect 10148 25540 10154 25542
rect 9846 25520 10154 25540
rect 10428 25158 10456 25842
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 9846 24508 10154 24528
rect 9846 24506 9852 24508
rect 9908 24506 9932 24508
rect 9988 24506 10012 24508
rect 10068 24506 10092 24508
rect 10148 24506 10154 24508
rect 9908 24454 9910 24506
rect 10090 24454 10092 24506
rect 9846 24452 9852 24454
rect 9908 24452 9932 24454
rect 9988 24452 10012 24454
rect 10068 24452 10092 24454
rect 10148 24452 10154 24454
rect 9846 24432 10154 24452
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7668 22234 7696 22578
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7852 21962 7880 23462
rect 8220 23050 8248 23666
rect 9846 23420 10154 23440
rect 9846 23418 9852 23420
rect 9908 23418 9932 23420
rect 9988 23418 10012 23420
rect 10068 23418 10092 23420
rect 10148 23418 10154 23420
rect 9908 23366 9910 23418
rect 10090 23366 10092 23418
rect 9846 23364 9852 23366
rect 9908 23364 9932 23366
rect 9988 23364 10012 23366
rect 10068 23364 10092 23366
rect 10148 23364 10154 23366
rect 9846 23344 10154 23364
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 8208 23044 8260 23050
rect 8208 22986 8260 22992
rect 8220 22094 8248 22986
rect 8312 22778 8340 23054
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8404 22710 8432 22918
rect 9140 22710 9168 23258
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 8128 22066 8248 22094
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 8128 21894 8156 22066
rect 8312 22030 8340 22510
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8128 20942 8156 21830
rect 8312 21554 8340 21966
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 8312 20942 8340 21490
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7668 20534 7696 20742
rect 7656 20528 7708 20534
rect 7656 20470 7708 20476
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7852 20058 7880 20402
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7248 17836 7328 17864
rect 7196 17818 7248 17824
rect 6644 17478 6696 17484
rect 6748 17496 6868 17524
rect 6656 17270 6684 17478
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6748 16250 6776 17496
rect 6880 17436 7188 17456
rect 6880 17434 6886 17436
rect 6942 17434 6966 17436
rect 7022 17434 7046 17436
rect 7102 17434 7126 17436
rect 7182 17434 7188 17436
rect 6942 17382 6944 17434
rect 7124 17382 7126 17434
rect 6880 17380 6886 17382
rect 6942 17380 6966 17382
rect 7022 17380 7046 17382
rect 7102 17380 7126 17382
rect 7182 17380 7188 17382
rect 6880 17360 7188 17380
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 7024 16794 7052 16934
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 7024 16658 7052 16730
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6880 16348 7188 16368
rect 6880 16346 6886 16348
rect 6942 16346 6966 16348
rect 7022 16346 7046 16348
rect 7102 16346 7126 16348
rect 7182 16346 7188 16348
rect 6942 16294 6944 16346
rect 7124 16294 7126 16346
rect 6880 16292 6886 16294
rect 6942 16292 6966 16294
rect 7022 16292 7046 16294
rect 7102 16292 7126 16294
rect 7182 16292 7188 16294
rect 6880 16272 7188 16292
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 7300 16182 7328 17836
rect 7484 17836 7604 17864
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7392 17134 7420 17546
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7392 16454 7420 17070
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6564 15570 6592 15846
rect 7300 15570 7328 16118
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 6564 15162 6592 15506
rect 7392 15434 7420 16390
rect 7484 15473 7512 17836
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7576 16590 7604 17682
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7470 15464 7526 15473
rect 7380 15428 7432 15434
rect 7470 15399 7526 15408
rect 7380 15370 7432 15376
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6288 10606 6316 11154
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 6288 10130 6316 10542
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5552 9654 5580 10066
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4540 8566 4568 8842
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3915 8188 4223 8208
rect 3915 8186 3921 8188
rect 3977 8186 4001 8188
rect 4057 8186 4081 8188
rect 4137 8186 4161 8188
rect 4217 8186 4223 8188
rect 3977 8134 3979 8186
rect 4159 8134 4161 8186
rect 3915 8132 3921 8134
rect 3977 8132 4001 8134
rect 4057 8132 4081 8134
rect 4137 8132 4161 8134
rect 4217 8132 4223 8134
rect 3915 8112 4223 8132
rect 3915 7100 4223 7120
rect 3915 7098 3921 7100
rect 3977 7098 4001 7100
rect 4057 7098 4081 7100
rect 4137 7098 4161 7100
rect 4217 7098 4223 7100
rect 3977 7046 3979 7098
rect 4159 7046 4161 7098
rect 3915 7044 3921 7046
rect 3977 7044 4001 7046
rect 4057 7044 4081 7046
rect 4137 7044 4161 7046
rect 4217 7044 4223 7046
rect 3915 7024 4223 7044
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 3915 6012 4223 6032
rect 3915 6010 3921 6012
rect 3977 6010 4001 6012
rect 4057 6010 4081 6012
rect 4137 6010 4161 6012
rect 4217 6010 4223 6012
rect 3977 5958 3979 6010
rect 4159 5958 4161 6010
rect 3915 5956 3921 5958
rect 3977 5956 4001 5958
rect 4057 5956 4081 5958
rect 4137 5956 4161 5958
rect 4217 5956 4223 5958
rect 3915 5936 4223 5956
rect 4540 5778 4568 6054
rect 5000 5914 5028 8842
rect 5276 8634 5304 9454
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5276 6322 5304 8570
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5552 6254 5580 9590
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 5552 5710 5580 6190
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5092 5370 5120 5646
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5448 5160 5500 5166
rect 5552 5114 5580 5510
rect 5500 5108 5580 5114
rect 5448 5102 5580 5108
rect 5356 5092 5408 5098
rect 5460 5086 5580 5102
rect 5356 5034 5408 5040
rect 3915 4924 4223 4944
rect 3915 4922 3921 4924
rect 3977 4922 4001 4924
rect 4057 4922 4081 4924
rect 4137 4922 4161 4924
rect 4217 4922 4223 4924
rect 3977 4870 3979 4922
rect 4159 4870 4161 4922
rect 3915 4868 3921 4870
rect 3977 4868 4001 4870
rect 4057 4868 4081 4870
rect 4137 4868 4161 4870
rect 4217 4868 4223 4870
rect 3915 4848 4223 4868
rect 5368 4622 5396 5034
rect 6380 5030 6408 9862
rect 6656 9654 6684 10066
rect 6748 9654 6776 15302
rect 6880 15260 7188 15280
rect 6880 15258 6886 15260
rect 6942 15258 6966 15260
rect 7022 15258 7046 15260
rect 7102 15258 7126 15260
rect 7182 15258 7188 15260
rect 6942 15206 6944 15258
rect 7124 15206 7126 15258
rect 6880 15204 6886 15206
rect 6942 15204 6966 15206
rect 7022 15204 7046 15206
rect 7102 15204 7126 15206
rect 7182 15204 7188 15206
rect 6880 15184 7188 15204
rect 7392 15026 7420 15370
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 6932 14550 6960 14962
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 6880 14172 7188 14192
rect 6880 14170 6886 14172
rect 6942 14170 6966 14172
rect 7022 14170 7046 14172
rect 7102 14170 7126 14172
rect 7182 14170 7188 14172
rect 6942 14118 6944 14170
rect 7124 14118 7126 14170
rect 6880 14116 6886 14118
rect 6942 14116 6966 14118
rect 7022 14116 7046 14118
rect 7102 14116 7126 14118
rect 7182 14116 7188 14118
rect 6880 14096 7188 14116
rect 6880 13084 7188 13104
rect 6880 13082 6886 13084
rect 6942 13082 6966 13084
rect 7022 13082 7046 13084
rect 7102 13082 7126 13084
rect 7182 13082 7188 13084
rect 6942 13030 6944 13082
rect 7124 13030 7126 13082
rect 6880 13028 6886 13030
rect 6942 13028 6966 13030
rect 7022 13028 7046 13030
rect 7102 13028 7126 13030
rect 7182 13028 7188 13030
rect 6880 13008 7188 13028
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 6880 11996 7188 12016
rect 6880 11994 6886 11996
rect 6942 11994 6966 11996
rect 7022 11994 7046 11996
rect 7102 11994 7126 11996
rect 7182 11994 7188 11996
rect 6942 11942 6944 11994
rect 7124 11942 7126 11994
rect 6880 11940 6886 11942
rect 6942 11940 6966 11942
rect 7022 11940 7046 11942
rect 7102 11940 7126 11942
rect 7182 11940 7188 11942
rect 6880 11920 7188 11940
rect 7300 11898 7328 12106
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7116 11558 7144 11766
rect 7576 11762 7604 16526
rect 7668 15638 7696 18158
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7668 14890 7696 15574
rect 7760 15026 7788 17546
rect 7852 16182 7880 19994
rect 8128 19854 8156 20878
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8220 17678 8248 18362
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 7840 16176 7892 16182
rect 7840 16118 7892 16124
rect 8036 16114 8064 16934
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 8036 15570 8064 16050
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8128 15434 8156 16118
rect 8220 15706 8248 17138
rect 8312 16794 8340 20878
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8404 17202 8432 20538
rect 8496 20330 8524 21490
rect 8588 20602 8616 21830
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 9048 20466 9076 22374
rect 9140 22030 9168 22646
rect 9324 22438 9352 22986
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9846 22332 10154 22352
rect 9846 22330 9852 22332
rect 9908 22330 9932 22332
rect 9988 22330 10012 22332
rect 10068 22330 10092 22332
rect 10148 22330 10154 22332
rect 9908 22278 9910 22330
rect 10090 22278 10092 22330
rect 9846 22276 9852 22278
rect 9908 22276 9932 22278
rect 9988 22276 10012 22278
rect 10068 22276 10092 22278
rect 10148 22276 10154 22278
rect 9846 22256 10154 22276
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9588 21956 9640 21962
rect 9588 21898 9640 21904
rect 9600 21350 9628 21898
rect 10244 21554 10272 23054
rect 10428 22094 10456 25094
rect 10520 24070 10548 34546
rect 10612 31346 10640 35634
rect 10796 33130 10824 38984
rect 10968 38820 11020 38826
rect 10968 38762 11020 38768
rect 10876 37936 10928 37942
rect 10876 37878 10928 37884
rect 10888 37398 10916 37878
rect 10980 37806 11008 38762
rect 11072 38486 11100 39034
rect 11060 38480 11112 38486
rect 11060 38422 11112 38428
rect 11612 38344 11664 38350
rect 11716 38332 11744 39374
rect 11808 38894 11836 39374
rect 12084 39098 12112 39986
rect 12268 39574 12296 43794
rect 12440 43716 12492 43722
rect 12440 43658 12492 43664
rect 12452 43450 12480 43658
rect 12532 43648 12584 43654
rect 12532 43590 12584 43596
rect 13268 43648 13320 43654
rect 13268 43590 13320 43596
rect 12440 43444 12492 43450
rect 12440 43386 12492 43392
rect 12544 43178 12572 43590
rect 12811 43548 13119 43568
rect 12811 43546 12817 43548
rect 12873 43546 12897 43548
rect 12953 43546 12977 43548
rect 13033 43546 13057 43548
rect 13113 43546 13119 43548
rect 12873 43494 12875 43546
rect 13055 43494 13057 43546
rect 12811 43492 12817 43494
rect 12873 43492 12897 43494
rect 12953 43492 12977 43494
rect 13033 43492 13057 43494
rect 13113 43492 13119 43494
rect 12811 43472 13119 43492
rect 12532 43172 12584 43178
rect 12532 43114 12584 43120
rect 12440 42696 12492 42702
rect 12440 42638 12492 42644
rect 12256 39568 12308 39574
rect 12256 39510 12308 39516
rect 12072 39092 12124 39098
rect 12072 39034 12124 39040
rect 12268 38962 12296 39510
rect 12452 39030 12480 42638
rect 12811 42460 13119 42480
rect 12811 42458 12817 42460
rect 12873 42458 12897 42460
rect 12953 42458 12977 42460
rect 13033 42458 13057 42460
rect 13113 42458 13119 42460
rect 12873 42406 12875 42458
rect 13055 42406 13057 42458
rect 12811 42404 12817 42406
rect 12873 42404 12897 42406
rect 12953 42404 12977 42406
rect 13033 42404 13057 42406
rect 13113 42404 13119 42406
rect 12811 42384 13119 42404
rect 12811 41372 13119 41392
rect 12811 41370 12817 41372
rect 12873 41370 12897 41372
rect 12953 41370 12977 41372
rect 13033 41370 13057 41372
rect 13113 41370 13119 41372
rect 12873 41318 12875 41370
rect 13055 41318 13057 41370
rect 12811 41316 12817 41318
rect 12873 41316 12897 41318
rect 12953 41316 12977 41318
rect 13033 41316 13057 41318
rect 13113 41316 13119 41318
rect 12811 41296 13119 41316
rect 12624 40520 12676 40526
rect 12624 40462 12676 40468
rect 12532 40044 12584 40050
rect 12532 39986 12584 39992
rect 12544 39506 12572 39986
rect 12636 39642 12664 40462
rect 12716 40384 12768 40390
rect 12716 40326 12768 40332
rect 12728 40118 12756 40326
rect 12811 40284 13119 40304
rect 12811 40282 12817 40284
rect 12873 40282 12897 40284
rect 12953 40282 12977 40284
rect 13033 40282 13057 40284
rect 13113 40282 13119 40284
rect 12873 40230 12875 40282
rect 13055 40230 13057 40282
rect 12811 40228 12817 40230
rect 12873 40228 12897 40230
rect 12953 40228 12977 40230
rect 13033 40228 13057 40230
rect 13113 40228 13119 40230
rect 12811 40208 13119 40228
rect 12716 40112 12768 40118
rect 12716 40054 12768 40060
rect 12624 39636 12676 39642
rect 12624 39578 12676 39584
rect 12532 39500 12584 39506
rect 12532 39442 12584 39448
rect 12440 39024 12492 39030
rect 12440 38966 12492 38972
rect 12256 38956 12308 38962
rect 12256 38898 12308 38904
rect 11796 38888 11848 38894
rect 11796 38830 11848 38836
rect 11808 38418 11836 38830
rect 11796 38412 11848 38418
rect 11796 38354 11848 38360
rect 12268 38350 12296 38898
rect 12452 38434 12480 38966
rect 12544 38554 12572 39442
rect 13176 39296 13228 39302
rect 13176 39238 13228 39244
rect 12811 39196 13119 39216
rect 12811 39194 12817 39196
rect 12873 39194 12897 39196
rect 12953 39194 12977 39196
rect 13033 39194 13057 39196
rect 13113 39194 13119 39196
rect 12873 39142 12875 39194
rect 13055 39142 13057 39194
rect 12811 39140 12817 39142
rect 12873 39140 12897 39142
rect 12953 39140 12977 39142
rect 13033 39140 13057 39142
rect 13113 39140 13119 39142
rect 12811 39120 13119 39140
rect 13188 38962 13216 39238
rect 13176 38956 13228 38962
rect 13176 38898 13228 38904
rect 12532 38548 12584 38554
rect 12532 38490 12584 38496
rect 12452 38406 12572 38434
rect 12544 38350 12572 38406
rect 11664 38304 11744 38332
rect 12256 38344 12308 38350
rect 11612 38286 11664 38292
rect 12256 38286 12308 38292
rect 12532 38344 12584 38350
rect 12532 38286 12584 38292
rect 12256 38208 12308 38214
rect 12256 38150 12308 38156
rect 11796 37868 11848 37874
rect 11796 37810 11848 37816
rect 10968 37800 11020 37806
rect 10968 37742 11020 37748
rect 10876 37392 10928 37398
rect 10876 37334 10928 37340
rect 10980 36174 11008 37742
rect 11808 37466 11836 37810
rect 11796 37460 11848 37466
rect 11796 37402 11848 37408
rect 12268 37262 12296 38150
rect 12544 38010 12572 38286
rect 12811 38108 13119 38128
rect 12811 38106 12817 38108
rect 12873 38106 12897 38108
rect 12953 38106 12977 38108
rect 13033 38106 13057 38108
rect 13113 38106 13119 38108
rect 12873 38054 12875 38106
rect 13055 38054 13057 38106
rect 12811 38052 12817 38054
rect 12873 38052 12897 38054
rect 12953 38052 12977 38054
rect 13033 38052 13057 38054
rect 13113 38052 13119 38054
rect 12811 38032 13119 38052
rect 12532 38004 12584 38010
rect 12532 37946 12584 37952
rect 11152 37256 11204 37262
rect 11152 37198 11204 37204
rect 12256 37256 12308 37262
rect 12256 37198 12308 37204
rect 10968 36168 11020 36174
rect 10968 36110 11020 36116
rect 10704 33114 10824 33130
rect 10692 33108 10824 33114
rect 10744 33102 10824 33108
rect 10692 33050 10744 33056
rect 10784 32836 10836 32842
rect 10784 32778 10836 32784
rect 10796 32502 10824 32778
rect 10784 32496 10836 32502
rect 10784 32438 10836 32444
rect 10796 31890 10824 32438
rect 10876 32224 10928 32230
rect 10876 32166 10928 32172
rect 10784 31884 10836 31890
rect 10784 31826 10836 31832
rect 10600 31340 10652 31346
rect 10600 31282 10652 31288
rect 10600 31204 10652 31210
rect 10600 31146 10652 31152
rect 10612 30734 10640 31146
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10612 30054 10640 30670
rect 10796 30258 10824 30738
rect 10784 30252 10836 30258
rect 10784 30194 10836 30200
rect 10600 30048 10652 30054
rect 10600 29990 10652 29996
rect 10888 28558 10916 32166
rect 10980 31482 11008 36110
rect 11164 35698 11192 37198
rect 12544 37194 12572 37946
rect 13280 37262 13308 43590
rect 13832 39982 13860 44338
rect 15776 44092 16084 44112
rect 15776 44090 15782 44092
rect 15838 44090 15862 44092
rect 15918 44090 15942 44092
rect 15998 44090 16022 44092
rect 16078 44090 16084 44092
rect 15838 44038 15840 44090
rect 16020 44038 16022 44090
rect 15776 44036 15782 44038
rect 15838 44036 15862 44038
rect 15918 44036 15942 44038
rect 15998 44036 16022 44038
rect 16078 44036 16084 44038
rect 15776 44016 16084 44036
rect 15776 43004 16084 43024
rect 15776 43002 15782 43004
rect 15838 43002 15862 43004
rect 15918 43002 15942 43004
rect 15998 43002 16022 43004
rect 16078 43002 16084 43004
rect 15838 42950 15840 43002
rect 16020 42950 16022 43002
rect 15776 42948 15782 42950
rect 15838 42948 15862 42950
rect 15918 42948 15942 42950
rect 15998 42948 16022 42950
rect 16078 42948 16084 42950
rect 15776 42928 16084 42948
rect 15776 41916 16084 41936
rect 15776 41914 15782 41916
rect 15838 41914 15862 41916
rect 15918 41914 15942 41916
rect 15998 41914 16022 41916
rect 16078 41914 16084 41916
rect 15838 41862 15840 41914
rect 16020 41862 16022 41914
rect 15776 41860 15782 41862
rect 15838 41860 15862 41862
rect 15918 41860 15942 41862
rect 15998 41860 16022 41862
rect 16078 41860 16084 41862
rect 15776 41840 16084 41860
rect 16672 41132 16724 41138
rect 16672 41074 16724 41080
rect 18144 41132 18196 41138
rect 18144 41074 18196 41080
rect 14464 41064 14516 41070
rect 14464 41006 14516 41012
rect 15384 41064 15436 41070
rect 15384 41006 15436 41012
rect 13820 39976 13872 39982
rect 13820 39918 13872 39924
rect 13832 39846 13860 39918
rect 14476 39846 14504 41006
rect 14740 40520 14792 40526
rect 14740 40462 14792 40468
rect 14648 40384 14700 40390
rect 14648 40326 14700 40332
rect 13820 39840 13872 39846
rect 13820 39782 13872 39788
rect 14464 39840 14516 39846
rect 14464 39782 14516 39788
rect 13452 39364 13504 39370
rect 13452 39306 13504 39312
rect 13360 38344 13412 38350
rect 13360 38286 13412 38292
rect 13372 37806 13400 38286
rect 13360 37800 13412 37806
rect 13360 37742 13412 37748
rect 13268 37256 13320 37262
rect 13268 37198 13320 37204
rect 12532 37188 12584 37194
rect 12532 37130 12584 37136
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 11152 35692 11204 35698
rect 11152 35634 11204 35640
rect 11796 34604 11848 34610
rect 11796 34546 11848 34552
rect 11520 34536 11572 34542
rect 11520 34478 11572 34484
rect 11532 33522 11560 34478
rect 11808 33862 11836 34546
rect 11980 34400 12032 34406
rect 11980 34342 12032 34348
rect 11796 33856 11848 33862
rect 11796 33798 11848 33804
rect 11808 33590 11836 33798
rect 11796 33584 11848 33590
rect 11796 33526 11848 33532
rect 11992 33522 12020 34342
rect 11520 33516 11572 33522
rect 11520 33458 11572 33464
rect 11980 33516 12032 33522
rect 11980 33458 12032 33464
rect 12256 33516 12308 33522
rect 12256 33458 12308 33464
rect 11532 33114 11560 33458
rect 11888 33312 11940 33318
rect 11888 33254 11940 33260
rect 11520 33108 11572 33114
rect 11520 33050 11572 33056
rect 11900 32570 11928 33254
rect 11888 32564 11940 32570
rect 11888 32506 11940 32512
rect 11900 32434 11928 32506
rect 11888 32428 11940 32434
rect 11888 32370 11940 32376
rect 11992 32298 12020 33458
rect 12072 33448 12124 33454
rect 12072 33390 12124 33396
rect 12084 32434 12112 33390
rect 12268 32434 12296 33458
rect 12072 32428 12124 32434
rect 12072 32370 12124 32376
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 11980 32292 12032 32298
rect 11980 32234 12032 32240
rect 12360 32230 12388 37062
rect 12811 37020 13119 37040
rect 12811 37018 12817 37020
rect 12873 37018 12897 37020
rect 12953 37018 12977 37020
rect 13033 37018 13057 37020
rect 13113 37018 13119 37020
rect 12873 36966 12875 37018
rect 13055 36966 13057 37018
rect 12811 36964 12817 36966
rect 12873 36964 12897 36966
rect 12953 36964 12977 36966
rect 13033 36964 13057 36966
rect 13113 36964 13119 36966
rect 12811 36944 13119 36964
rect 12716 36780 12768 36786
rect 12716 36722 12768 36728
rect 12728 34542 12756 36722
rect 12811 35932 13119 35952
rect 12811 35930 12817 35932
rect 12873 35930 12897 35932
rect 12953 35930 12977 35932
rect 13033 35930 13057 35932
rect 13113 35930 13119 35932
rect 12873 35878 12875 35930
rect 13055 35878 13057 35930
rect 12811 35876 12817 35878
rect 12873 35876 12897 35878
rect 12953 35876 12977 35878
rect 13033 35876 13057 35878
rect 13113 35876 13119 35878
rect 12811 35856 13119 35876
rect 12811 34844 13119 34864
rect 12811 34842 12817 34844
rect 12873 34842 12897 34844
rect 12953 34842 12977 34844
rect 13033 34842 13057 34844
rect 13113 34842 13119 34844
rect 12873 34790 12875 34842
rect 13055 34790 13057 34842
rect 12811 34788 12817 34790
rect 12873 34788 12897 34790
rect 12953 34788 12977 34790
rect 13033 34788 13057 34790
rect 13113 34788 13119 34790
rect 12811 34768 13119 34788
rect 12716 34536 12768 34542
rect 12716 34478 12768 34484
rect 12440 33380 12492 33386
rect 12440 33322 12492 33328
rect 12452 32366 12480 33322
rect 12624 32836 12676 32842
rect 12624 32778 12676 32784
rect 12440 32360 12492 32366
rect 12440 32302 12492 32308
rect 12348 32224 12400 32230
rect 12348 32166 12400 32172
rect 12452 31890 12480 32302
rect 12636 32026 12664 32778
rect 12728 32502 12756 34478
rect 13176 34400 13228 34406
rect 13176 34342 13228 34348
rect 12811 33756 13119 33776
rect 12811 33754 12817 33756
rect 12873 33754 12897 33756
rect 12953 33754 12977 33756
rect 13033 33754 13057 33756
rect 13113 33754 13119 33756
rect 12873 33702 12875 33754
rect 13055 33702 13057 33754
rect 12811 33700 12817 33702
rect 12873 33700 12897 33702
rect 12953 33700 12977 33702
rect 13033 33700 13057 33702
rect 13113 33700 13119 33702
rect 12811 33680 13119 33700
rect 13188 33590 13216 34342
rect 13360 33992 13412 33998
rect 13360 33934 13412 33940
rect 13176 33584 13228 33590
rect 13176 33526 13228 33532
rect 13188 32978 13216 33526
rect 13176 32972 13228 32978
rect 13176 32914 13228 32920
rect 12811 32668 13119 32688
rect 12811 32666 12817 32668
rect 12873 32666 12897 32668
rect 12953 32666 12977 32668
rect 13033 32666 13057 32668
rect 13113 32666 13119 32668
rect 12873 32614 12875 32666
rect 13055 32614 13057 32666
rect 12811 32612 12817 32614
rect 12873 32612 12897 32614
rect 12953 32612 12977 32614
rect 13033 32612 13057 32614
rect 13113 32612 13119 32614
rect 12811 32592 13119 32612
rect 12716 32496 12768 32502
rect 12716 32438 12768 32444
rect 13188 32298 13216 32914
rect 13372 32910 13400 33934
rect 13360 32904 13412 32910
rect 13360 32846 13412 32852
rect 13176 32292 13228 32298
rect 13176 32234 13228 32240
rect 12624 32020 12676 32026
rect 12624 31962 12676 31968
rect 12440 31884 12492 31890
rect 12440 31826 12492 31832
rect 11796 31816 11848 31822
rect 11796 31758 11848 31764
rect 12452 31770 12480 31826
rect 11152 31748 11204 31754
rect 11152 31690 11204 31696
rect 10968 31476 11020 31482
rect 10968 31418 11020 31424
rect 11164 31346 11192 31690
rect 11152 31340 11204 31346
rect 11152 31282 11204 31288
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 10980 30666 11008 31078
rect 10968 30660 11020 30666
rect 10968 30602 11020 30608
rect 11336 30184 11388 30190
rect 11336 30126 11388 30132
rect 11348 29646 11376 30126
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 11348 27470 11376 29582
rect 11336 27464 11388 27470
rect 11336 27406 11388 27412
rect 11612 27464 11664 27470
rect 11612 27406 11664 27412
rect 10692 26240 10744 26246
rect 10692 26182 10744 26188
rect 10704 25906 10732 26182
rect 11348 25974 11376 27406
rect 11624 27130 11652 27406
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11704 26852 11756 26858
rect 11704 26794 11756 26800
rect 11716 26382 11744 26794
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 11336 25968 11388 25974
rect 11336 25910 11388 25916
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 11612 25832 11664 25838
rect 11612 25774 11664 25780
rect 11624 25430 11652 25774
rect 11612 25424 11664 25430
rect 11612 25366 11664 25372
rect 11520 25220 11572 25226
rect 11520 25162 11572 25168
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 11336 25152 11388 25158
rect 11336 25094 11388 25100
rect 11164 24886 11192 25094
rect 11152 24880 11204 24886
rect 11152 24822 11204 24828
rect 10508 24064 10560 24070
rect 10508 24006 10560 24012
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10520 22642 10548 22918
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 10428 22066 10640 22094
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9600 20874 9628 21286
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9508 20534 9536 20742
rect 9496 20528 9548 20534
rect 9496 20470 9548 20476
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8588 17202 8616 20198
rect 9508 19854 9536 20470
rect 9692 20262 9720 21422
rect 9846 21244 10154 21264
rect 9846 21242 9852 21244
rect 9908 21242 9932 21244
rect 9988 21242 10012 21244
rect 10068 21242 10092 21244
rect 10148 21242 10154 21244
rect 9908 21190 9910 21242
rect 10090 21190 10092 21242
rect 9846 21188 9852 21190
rect 9908 21188 9932 21190
rect 9988 21188 10012 21190
rect 10068 21188 10092 21190
rect 10148 21188 10154 21190
rect 9846 21168 10154 21188
rect 10244 20602 10272 21490
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8404 15994 8432 17138
rect 8588 16250 8616 17138
rect 8772 16590 8800 17138
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8312 15966 8432 15994
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8312 15638 8340 15966
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8404 15502 8432 15846
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7380 11756 7432 11762
rect 7564 11756 7616 11762
rect 7380 11698 7432 11704
rect 7484 11716 7564 11744
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7392 11354 7420 11698
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7392 11082 7420 11154
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 6880 10908 7188 10928
rect 6880 10906 6886 10908
rect 6942 10906 6966 10908
rect 7022 10906 7046 10908
rect 7102 10906 7126 10908
rect 7182 10906 7188 10908
rect 6942 10854 6944 10906
rect 7124 10854 7126 10906
rect 6880 10852 6886 10854
rect 6942 10852 6966 10854
rect 7022 10852 7046 10854
rect 7102 10852 7126 10854
rect 7182 10852 7188 10854
rect 6880 10832 7188 10852
rect 7300 10538 7328 11018
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7024 10266 7052 10474
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7012 10056 7064 10062
rect 7010 10024 7012 10033
rect 7064 10024 7066 10033
rect 7300 10010 7328 10134
rect 7010 9959 7066 9968
rect 7291 9982 7328 10010
rect 6880 9820 7188 9840
rect 6880 9818 6886 9820
rect 6942 9818 6966 9820
rect 7022 9818 7046 9820
rect 7102 9818 7126 9820
rect 7182 9818 7188 9820
rect 6942 9766 6944 9818
rect 7124 9766 7126 9818
rect 6880 9764 6886 9766
rect 6942 9764 6966 9766
rect 7022 9764 7046 9766
rect 7102 9764 7126 9766
rect 7182 9764 7188 9766
rect 6880 9744 7188 9764
rect 7102 9688 7158 9697
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6736 9648 6788 9654
rect 7291 9674 7319 9982
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7291 9646 7328 9674
rect 7102 9623 7158 9632
rect 6736 9590 6788 9596
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 7116 8922 7144 9623
rect 7300 9586 7328 9646
rect 7392 9586 7420 9862
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 6564 6390 6592 8910
rect 7116 8894 7328 8922
rect 6880 8732 7188 8752
rect 6880 8730 6886 8732
rect 6942 8730 6966 8732
rect 7022 8730 7046 8732
rect 7102 8730 7126 8732
rect 7182 8730 7188 8732
rect 6942 8678 6944 8730
rect 7124 8678 7126 8730
rect 6880 8676 6886 8678
rect 6942 8676 6966 8678
rect 7022 8676 7046 8678
rect 7102 8676 7126 8678
rect 7182 8676 7188 8678
rect 6880 8656 7188 8676
rect 6880 7644 7188 7664
rect 6880 7642 6886 7644
rect 6942 7642 6966 7644
rect 7022 7642 7046 7644
rect 7102 7642 7126 7644
rect 7182 7642 7188 7644
rect 6942 7590 6944 7642
rect 7124 7590 7126 7642
rect 6880 7588 6886 7590
rect 6942 7588 6966 7590
rect 7022 7588 7046 7590
rect 7102 7588 7126 7590
rect 7182 7588 7188 7590
rect 6880 7568 7188 7588
rect 6880 6556 7188 6576
rect 6880 6554 6886 6556
rect 6942 6554 6966 6556
rect 7022 6554 7046 6556
rect 7102 6554 7126 6556
rect 7182 6554 7188 6556
rect 6942 6502 6944 6554
rect 7124 6502 7126 6554
rect 6880 6500 6886 6502
rect 6942 6500 6966 6502
rect 7022 6500 7046 6502
rect 7102 6500 7126 6502
rect 7182 6500 7188 6502
rect 6880 6480 7188 6500
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 5552 4690 5580 4966
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 6564 4486 6592 6326
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6748 5914 6776 6258
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6656 5710 6684 5782
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5234 6684 5646
rect 7300 5642 7328 8894
rect 7392 8498 7420 9522
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7484 6798 7512 11716
rect 7564 11698 7616 11704
rect 7668 11218 7696 14826
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7760 11098 7788 14962
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7668 11070 7788 11098
rect 7668 10742 7696 11070
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7760 10742 7788 10950
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 10130 7696 10406
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7760 9994 7788 10678
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7760 9654 7788 9930
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7472 6792 7524 6798
rect 7392 6752 7472 6780
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 6748 5302 6776 5578
rect 6880 5468 7188 5488
rect 6880 5466 6886 5468
rect 6942 5466 6966 5468
rect 7022 5466 7046 5468
rect 7102 5466 7126 5468
rect 7182 5466 7188 5468
rect 6942 5414 6944 5466
rect 7124 5414 7126 5466
rect 6880 5412 6886 5414
rect 6942 5412 6966 5414
rect 7022 5412 7046 5414
rect 7102 5412 7126 5414
rect 7182 5412 7188 5414
rect 6880 5392 7188 5412
rect 7392 5302 7420 6752
rect 7472 6734 7524 6740
rect 7576 6322 7604 9522
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7668 6322 7696 9386
rect 7852 8974 7880 14486
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 11150 7972 11494
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7944 10810 7972 11086
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8036 9110 8064 11562
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8220 9738 8248 10610
rect 8404 10062 8432 15030
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8588 12918 8616 14962
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8588 12442 8616 12854
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8680 12170 8708 12582
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8680 11830 8708 12106
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11150 8708 11494
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8392 10056 8444 10062
rect 8772 10033 8800 16526
rect 8956 14618 8984 16934
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 9140 14414 9168 14758
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 12238 8984 14214
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8864 11218 8892 12174
rect 9048 11762 9076 12310
rect 9232 12238 9260 14894
rect 9324 14006 9352 16594
rect 9508 14958 9536 19654
rect 9692 19378 9720 20198
rect 9846 20156 10154 20176
rect 9846 20154 9852 20156
rect 9908 20154 9932 20156
rect 9988 20154 10012 20156
rect 10068 20154 10092 20156
rect 10148 20154 10154 20156
rect 9908 20102 9910 20154
rect 10090 20102 10092 20154
rect 9846 20100 9852 20102
rect 9908 20100 9932 20102
rect 9988 20100 10012 20102
rect 10068 20100 10092 20102
rect 10148 20100 10154 20102
rect 9846 20080 10154 20100
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9692 17678 9720 17750
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16522 9720 16934
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9600 14482 9628 15846
rect 9692 15094 9720 16118
rect 9784 16114 9812 19382
rect 9846 19068 10154 19088
rect 9846 19066 9852 19068
rect 9908 19066 9932 19068
rect 9988 19066 10012 19068
rect 10068 19066 10092 19068
rect 10148 19066 10154 19068
rect 9908 19014 9910 19066
rect 10090 19014 10092 19066
rect 9846 19012 9852 19014
rect 9908 19012 9932 19014
rect 9988 19012 10012 19014
rect 10068 19012 10092 19014
rect 10148 19012 10154 19014
rect 9846 18992 10154 19012
rect 9846 17980 10154 18000
rect 9846 17978 9852 17980
rect 9908 17978 9932 17980
rect 9988 17978 10012 17980
rect 10068 17978 10092 17980
rect 10148 17978 10154 17980
rect 9908 17926 9910 17978
rect 10090 17926 10092 17978
rect 9846 17924 9852 17926
rect 9908 17924 9932 17926
rect 9988 17924 10012 17926
rect 10068 17924 10092 17926
rect 10148 17924 10154 17926
rect 9846 17904 10154 17924
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9876 17202 9904 17478
rect 10244 17202 10272 20198
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 9846 16892 10154 16912
rect 9846 16890 9852 16892
rect 9908 16890 9932 16892
rect 9988 16890 10012 16892
rect 10068 16890 10092 16892
rect 10148 16890 10154 16892
rect 9908 16838 9910 16890
rect 10090 16838 10092 16890
rect 9846 16836 9852 16838
rect 9908 16836 9932 16838
rect 9988 16836 10012 16838
rect 10068 16836 10092 16838
rect 10148 16836 10154 16838
rect 9846 16816 10154 16836
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16114 10180 16526
rect 10244 16182 10272 17138
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9784 15026 9812 16050
rect 9846 15804 10154 15824
rect 9846 15802 9852 15804
rect 9908 15802 9932 15804
rect 9988 15802 10012 15804
rect 10068 15802 10092 15804
rect 10148 15802 10154 15804
rect 9908 15750 9910 15802
rect 10090 15750 10092 15802
rect 9846 15748 9852 15750
rect 9908 15748 9932 15750
rect 9988 15748 10012 15750
rect 10068 15748 10092 15750
rect 10148 15748 10154 15750
rect 9846 15728 10154 15748
rect 10244 15162 10272 16118
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10336 15094 10364 15302
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10244 14890 10272 14962
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 9846 14716 10154 14736
rect 9846 14714 9852 14716
rect 9908 14714 9932 14716
rect 9988 14714 10012 14716
rect 10068 14714 10092 14716
rect 10148 14714 10154 14716
rect 9908 14662 9910 14714
rect 10090 14662 10092 14714
rect 9846 14660 9852 14662
rect 9908 14660 9932 14662
rect 9988 14660 10012 14662
rect 10068 14660 10092 14662
rect 10148 14660 10154 14662
rect 9846 14640 10154 14660
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9600 12306 9628 12582
rect 9692 12322 9720 14214
rect 9876 14006 9904 14282
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9876 13818 9904 13942
rect 9784 13790 9904 13818
rect 9784 12918 9812 13790
rect 9846 13628 10154 13648
rect 9846 13626 9852 13628
rect 9908 13626 9932 13628
rect 9988 13626 10012 13628
rect 10068 13626 10092 13628
rect 10148 13626 10154 13628
rect 9908 13574 9910 13626
rect 10090 13574 10092 13626
rect 9846 13572 9852 13574
rect 9908 13572 9932 13574
rect 9988 13572 10012 13574
rect 10068 13572 10092 13574
rect 10148 13572 10154 13574
rect 9846 13552 10154 13572
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 12434 9812 12582
rect 9846 12540 10154 12560
rect 9846 12538 9852 12540
rect 9908 12538 9932 12540
rect 9988 12538 10012 12540
rect 10068 12538 10092 12540
rect 10148 12538 10154 12540
rect 9908 12486 9910 12538
rect 10090 12486 10092 12538
rect 9846 12484 9852 12486
rect 9908 12484 9932 12486
rect 9988 12484 10012 12486
rect 10068 12484 10092 12486
rect 10148 12484 10154 12486
rect 9846 12464 10154 12484
rect 10244 12434 10272 14826
rect 10336 12850 10364 15030
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 9784 12406 9904 12434
rect 9588 12300 9640 12306
rect 9692 12294 9812 12322
rect 9588 12242 9640 12248
rect 9784 12238 9812 12294
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8392 9998 8444 10004
rect 8758 10024 8814 10033
rect 8220 9710 8340 9738
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 8036 8514 8064 9046
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 7840 8492 7892 8498
rect 8036 8486 8156 8514
rect 7840 8434 7892 8440
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7886 7788 8230
rect 7852 7886 7880 8434
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7760 6458 7788 7822
rect 7840 6792 7892 6798
rect 7944 6780 7972 8298
rect 8036 8090 8064 8366
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8128 6866 8156 8486
rect 8220 7954 8248 8910
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7892 6752 7972 6780
rect 7840 6734 7892 6740
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 8128 6338 8156 6802
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 8036 6310 8156 6338
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6656 4758 6684 5170
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 7392 4622 7420 5238
rect 7484 5234 7512 6054
rect 7576 5710 7604 6258
rect 7668 5778 7696 6258
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 5736 4146 5764 4422
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 3915 3836 4223 3856
rect 3915 3834 3921 3836
rect 3977 3834 4001 3836
rect 4057 3834 4081 3836
rect 4137 3834 4161 3836
rect 4217 3834 4223 3836
rect 3977 3782 3979 3834
rect 4159 3782 4161 3834
rect 3915 3780 3921 3782
rect 3977 3780 4001 3782
rect 4057 3780 4081 3782
rect 4137 3780 4161 3782
rect 4217 3780 4223 3782
rect 3915 3760 4223 3780
rect 6104 3602 6132 4014
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6196 3534 6224 4422
rect 6564 4146 6592 4422
rect 6656 4282 6684 4558
rect 6880 4380 7188 4400
rect 6880 4378 6886 4380
rect 6942 4378 6966 4380
rect 7022 4378 7046 4380
rect 7102 4378 7126 4380
rect 7182 4378 7188 4380
rect 6942 4326 6944 4378
rect 7124 4326 7126 4378
rect 6880 4324 6886 4326
rect 6942 4324 6966 4326
rect 7022 4324 7046 4326
rect 7102 4324 7126 4326
rect 7182 4324 7188 4326
rect 6880 4304 7188 4324
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 7484 3738 7512 4694
rect 7576 4146 7604 4966
rect 7668 4826 7696 5714
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7760 5234 7788 5578
rect 8036 5302 8064 6310
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 5574 8156 6190
rect 8312 5710 8340 9710
rect 8404 7562 8432 9998
rect 8758 9959 8814 9968
rect 8864 9586 8892 11154
rect 9232 10674 9260 11766
rect 9324 11014 9352 12106
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10742 9352 10950
rect 9600 10810 9628 11698
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9692 10674 9720 12038
rect 9784 10742 9812 12174
rect 9876 11830 9904 12406
rect 10152 12406 10272 12434
rect 10152 12238 10180 12406
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9968 11762 9996 11834
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 10152 11626 10180 12174
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 9846 11452 10154 11472
rect 9846 11450 9852 11452
rect 9908 11450 9932 11452
rect 9988 11450 10012 11452
rect 10068 11450 10092 11452
rect 10148 11450 10154 11452
rect 9908 11398 9910 11450
rect 10090 11398 10092 11450
rect 9846 11396 9852 11398
rect 9908 11396 9932 11398
rect 9988 11396 10012 11398
rect 10068 11396 10092 11398
rect 10148 11396 10154 11398
rect 9846 11376 10154 11396
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8404 7546 8524 7562
rect 8404 7540 8536 7546
rect 8404 7534 8484 7540
rect 8484 7482 8536 7488
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 7002 8432 7346
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8496 6798 8524 7482
rect 8864 7478 8892 9522
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8864 6866 8892 7414
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 9232 5846 9260 10610
rect 10244 10606 10272 11766
rect 10336 11694 10364 12038
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 11354 10364 11630
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10336 10674 10364 11290
rect 10428 10810 10456 15982
rect 10520 12170 10548 17750
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10520 10470 10548 11834
rect 10612 10606 10640 22066
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 10704 21690 10732 22034
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10704 19990 10732 21626
rect 10980 21486 11008 21830
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 11256 21010 11284 22510
rect 11348 22094 11376 25094
rect 11532 22642 11560 25162
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11348 22066 11560 22094
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10796 20058 10824 20810
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10692 19984 10744 19990
rect 10692 19926 10744 19932
rect 10980 19854 11008 20198
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10704 16794 10732 17070
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10704 16114 10732 16730
rect 10980 16250 11008 17614
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11164 17066 11192 17546
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10704 14822 10732 16050
rect 10980 15706 11008 16186
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10888 15162 10916 15370
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10704 14414 10732 14758
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 11164 11218 11192 17002
rect 11256 16794 11284 20946
rect 11348 20398 11376 21286
rect 11440 20602 11468 21966
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 11348 19922 11376 20334
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11256 16658 11284 16730
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11256 15570 11284 16594
rect 11348 15570 11376 19858
rect 11532 17882 11560 22066
rect 11624 20942 11652 22374
rect 11716 21350 11744 26318
rect 11808 25294 11836 31758
rect 12452 31742 12572 31770
rect 12544 29850 12572 31742
rect 12811 31580 13119 31600
rect 12811 31578 12817 31580
rect 12873 31578 12897 31580
rect 12953 31578 12977 31580
rect 13033 31578 13057 31580
rect 13113 31578 13119 31580
rect 12873 31526 12875 31578
rect 13055 31526 13057 31578
rect 12811 31524 12817 31526
rect 12873 31524 12897 31526
rect 12953 31524 12977 31526
rect 13033 31524 13057 31526
rect 13113 31524 13119 31526
rect 12811 31504 13119 31524
rect 13360 31136 13412 31142
rect 13360 31078 13412 31084
rect 13372 30734 13400 31078
rect 13360 30728 13412 30734
rect 13360 30670 13412 30676
rect 12811 30492 13119 30512
rect 12811 30490 12817 30492
rect 12873 30490 12897 30492
rect 12953 30490 12977 30492
rect 13033 30490 13057 30492
rect 13113 30490 13119 30492
rect 12873 30438 12875 30490
rect 13055 30438 13057 30490
rect 12811 30436 12817 30438
rect 12873 30436 12897 30438
rect 12953 30436 12977 30438
rect 13033 30436 13057 30438
rect 13113 30436 13119 30438
rect 12811 30416 13119 30436
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 12084 28762 12112 29514
rect 12072 28756 12124 28762
rect 12072 28698 12124 28704
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 11888 28076 11940 28082
rect 11888 28018 11940 28024
rect 11900 27402 11928 28018
rect 12360 27470 12388 28494
rect 12544 28218 12572 29786
rect 13360 29640 13412 29646
rect 13360 29582 13412 29588
rect 12811 29404 13119 29424
rect 12811 29402 12817 29404
rect 12873 29402 12897 29404
rect 12953 29402 12977 29404
rect 13033 29402 13057 29404
rect 13113 29402 13119 29404
rect 12873 29350 12875 29402
rect 13055 29350 13057 29402
rect 12811 29348 12817 29350
rect 12873 29348 12897 29350
rect 12953 29348 12977 29350
rect 13033 29348 13057 29350
rect 13113 29348 13119 29350
rect 12811 29328 13119 29348
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12440 28076 12492 28082
rect 12440 28018 12492 28024
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 11888 27396 11940 27402
rect 11888 27338 11940 27344
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11900 21554 11928 27338
rect 12256 27328 12308 27334
rect 12256 27270 12308 27276
rect 12268 26994 12296 27270
rect 12452 27130 12480 28018
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12532 27056 12584 27062
rect 12532 26998 12584 27004
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 12084 26586 12112 26930
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 12072 25424 12124 25430
rect 12072 25366 12124 25372
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11900 20534 11928 21490
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11532 14482 11560 17478
rect 11716 17134 11744 17614
rect 11808 17202 11836 17750
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11900 15366 11928 16458
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11716 15026 11744 15302
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11624 12238 11652 12718
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11624 11762 11652 12174
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11440 10810 11468 11290
rect 11532 11014 11560 11494
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 9846 10364 10154 10384
rect 9846 10362 9852 10364
rect 9908 10362 9932 10364
rect 9988 10362 10012 10364
rect 10068 10362 10092 10364
rect 10148 10362 10154 10364
rect 9908 10310 9910 10362
rect 10090 10310 10092 10362
rect 9846 10308 9852 10310
rect 9908 10308 9932 10310
rect 9988 10308 10012 10310
rect 10068 10308 10092 10310
rect 10148 10308 10154 10310
rect 9846 10288 10154 10308
rect 10520 9654 10548 10406
rect 11808 10266 11836 12106
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 9846 9276 10154 9296
rect 9846 9274 9852 9276
rect 9908 9274 9932 9276
rect 9988 9274 10012 9276
rect 10068 9274 10092 9276
rect 10148 9274 10154 9276
rect 9908 9222 9910 9274
rect 10090 9222 10092 9274
rect 9846 9220 9852 9222
rect 9908 9220 9932 9222
rect 9988 9220 10012 9222
rect 10068 9220 10092 9222
rect 10148 9220 10154 9222
rect 9846 9200 10154 9220
rect 10244 9178 10272 9522
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10428 8634 10456 8910
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10520 8430 10548 8978
rect 10704 8974 10732 9318
rect 11440 9178 11468 9998
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 9846 8188 10154 8208
rect 9846 8186 9852 8188
rect 9908 8186 9932 8188
rect 9988 8186 10012 8188
rect 10068 8186 10092 8188
rect 10148 8186 10154 8188
rect 9908 8134 9910 8186
rect 10090 8134 10092 8186
rect 9846 8132 9852 8134
rect 9908 8132 9932 8134
rect 9988 8132 10012 8134
rect 10068 8132 10092 8134
rect 10148 8132 10154 8134
rect 9846 8112 10154 8132
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 9846 7100 10154 7120
rect 9846 7098 9852 7100
rect 9908 7098 9932 7100
rect 9988 7098 10012 7100
rect 10068 7098 10092 7100
rect 10148 7098 10154 7100
rect 9908 7046 9910 7098
rect 10090 7046 10092 7098
rect 9846 7044 9852 7046
rect 9908 7044 9932 7046
rect 9988 7044 10012 7046
rect 10068 7044 10092 7046
rect 10148 7044 10154 7046
rect 9846 7024 10154 7044
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9508 5778 9536 6802
rect 10244 6798 10272 7142
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7760 4826 7788 5170
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 8128 4690 8156 5510
rect 8312 5370 8340 5646
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8312 4554 8340 5170
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8404 4622 8432 4966
rect 9508 4690 9536 5714
rect 9784 5710 9812 6598
rect 9846 6012 10154 6032
rect 9846 6010 9852 6012
rect 9908 6010 9932 6012
rect 9988 6010 10012 6012
rect 10068 6010 10092 6012
rect 10148 6010 10154 6012
rect 9908 5958 9910 6010
rect 10090 5958 10092 6010
rect 9846 5956 9852 5958
rect 9908 5956 9932 5958
rect 9988 5956 10012 5958
rect 10068 5956 10092 5958
rect 10148 5956 10154 5958
rect 9846 5936 10154 5956
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8312 4282 8340 4490
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 9508 4214 9536 4626
rect 9692 4622 9720 4966
rect 9846 4924 10154 4944
rect 9846 4922 9852 4924
rect 9908 4922 9932 4924
rect 9988 4922 10012 4924
rect 10068 4922 10092 4924
rect 10148 4922 10154 4924
rect 9908 4870 9910 4922
rect 10090 4870 10092 4922
rect 9846 4868 9852 4870
rect 9908 4868 9932 4870
rect 9988 4868 10012 4870
rect 10068 4868 10092 4870
rect 10148 4868 10154 4870
rect 9846 4848 10154 4868
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 10520 4282 10548 8366
rect 10704 8362 10732 8910
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10704 7410 10732 8298
rect 10980 8242 11008 8434
rect 10980 8214 11100 8242
rect 11072 7750 11100 8214
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 11072 7342 11100 7686
rect 11532 7546 11560 8910
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10888 5914 10916 7142
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10888 5234 10916 5850
rect 11072 5710 11100 7278
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 11072 5166 11100 5646
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9784 3738 9812 4082
rect 9846 3836 10154 3856
rect 9846 3834 9852 3836
rect 9908 3834 9932 3836
rect 9988 3834 10012 3836
rect 10068 3834 10092 3836
rect 10148 3834 10154 3836
rect 9908 3782 9910 3834
rect 10090 3782 10092 3834
rect 9846 3780 9852 3782
rect 9908 3780 9932 3782
rect 9988 3780 10012 3782
rect 10068 3780 10092 3782
rect 10148 3780 10154 3782
rect 9846 3760 10154 3780
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 11072 3534 11100 5102
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11164 3602 11192 4762
rect 11440 4690 11468 6802
rect 11624 6458 11652 9998
rect 11900 8974 11928 15302
rect 11992 15094 12020 24006
rect 12084 22094 12112 25366
rect 12268 25362 12296 26930
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 12452 26450 12480 26726
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12544 25294 12572 26998
rect 12636 26926 12664 28562
rect 13372 28558 13400 29582
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 12728 28218 12756 28494
rect 12811 28316 13119 28336
rect 12811 28314 12817 28316
rect 12873 28314 12897 28316
rect 12953 28314 12977 28316
rect 13033 28314 13057 28316
rect 13113 28314 13119 28316
rect 12873 28262 12875 28314
rect 13055 28262 13057 28314
rect 12811 28260 12817 28262
rect 12873 28260 12897 28262
rect 12953 28260 12977 28262
rect 13033 28260 13057 28262
rect 13113 28260 13119 28262
rect 12811 28240 13119 28260
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 13360 27668 13412 27674
rect 13360 27610 13412 27616
rect 12811 27228 13119 27248
rect 12811 27226 12817 27228
rect 12873 27226 12897 27228
rect 12953 27226 12977 27228
rect 13033 27226 13057 27228
rect 13113 27226 13119 27228
rect 12873 27174 12875 27226
rect 13055 27174 13057 27226
rect 12811 27172 12817 27174
rect 12873 27172 12897 27174
rect 12953 27172 12977 27174
rect 13033 27172 13057 27174
rect 13113 27172 13119 27174
rect 12811 27152 13119 27172
rect 13372 27062 13400 27610
rect 13360 27056 13412 27062
rect 13360 26998 13412 27004
rect 12624 26920 12676 26926
rect 12624 26862 12676 26868
rect 12636 26042 12664 26862
rect 13464 26858 13492 39306
rect 13832 39030 13860 39782
rect 14660 39438 14688 40326
rect 14752 39982 14780 40462
rect 15396 40118 15424 41006
rect 15476 40928 15528 40934
rect 15476 40870 15528 40876
rect 16120 40928 16172 40934
rect 16120 40870 16172 40876
rect 15488 40458 15516 40870
rect 15776 40828 16084 40848
rect 15776 40826 15782 40828
rect 15838 40826 15862 40828
rect 15918 40826 15942 40828
rect 15998 40826 16022 40828
rect 16078 40826 16084 40828
rect 15838 40774 15840 40826
rect 16020 40774 16022 40826
rect 15776 40772 15782 40774
rect 15838 40772 15862 40774
rect 15918 40772 15942 40774
rect 15998 40772 16022 40774
rect 16078 40772 16084 40774
rect 15776 40752 16084 40772
rect 16132 40526 16160 40870
rect 16120 40520 16172 40526
rect 16120 40462 16172 40468
rect 15476 40452 15528 40458
rect 15476 40394 15528 40400
rect 15384 40112 15436 40118
rect 15384 40054 15436 40060
rect 14740 39976 14792 39982
rect 14740 39918 14792 39924
rect 15108 39840 15160 39846
rect 15108 39782 15160 39788
rect 15120 39642 15148 39782
rect 15396 39642 15424 40054
rect 15568 40044 15620 40050
rect 15568 39986 15620 39992
rect 15108 39636 15160 39642
rect 15108 39578 15160 39584
rect 15384 39636 15436 39642
rect 15384 39578 15436 39584
rect 14648 39432 14700 39438
rect 14648 39374 14700 39380
rect 14188 39364 14240 39370
rect 14188 39306 14240 39312
rect 13820 39024 13872 39030
rect 13820 38966 13872 38972
rect 13832 38418 13860 38966
rect 14200 38962 14228 39306
rect 14660 39030 14688 39374
rect 14924 39296 14976 39302
rect 14924 39238 14976 39244
rect 14648 39024 14700 39030
rect 14648 38966 14700 38972
rect 14188 38956 14240 38962
rect 14188 38898 14240 38904
rect 14200 38758 14228 38898
rect 14188 38752 14240 38758
rect 14188 38694 14240 38700
rect 14372 38752 14424 38758
rect 14372 38694 14424 38700
rect 13820 38412 13872 38418
rect 13820 38354 13872 38360
rect 13832 37942 13860 38354
rect 13820 37936 13872 37942
rect 13820 37878 13872 37884
rect 13832 36922 13860 37878
rect 14200 37874 14228 38694
rect 14004 37868 14056 37874
rect 14004 37810 14056 37816
rect 14188 37868 14240 37874
rect 14188 37810 14240 37816
rect 13820 36916 13872 36922
rect 13820 36858 13872 36864
rect 13832 35630 13860 36858
rect 13820 35624 13872 35630
rect 13820 35566 13872 35572
rect 14016 33522 14044 37810
rect 14384 35086 14412 38694
rect 14936 36174 14964 39238
rect 15120 39098 15148 39578
rect 15200 39500 15252 39506
rect 15200 39442 15252 39448
rect 15108 39092 15160 39098
rect 15108 39034 15160 39040
rect 15212 38962 15240 39442
rect 15200 38956 15252 38962
rect 15200 38898 15252 38904
rect 15212 38554 15240 38898
rect 15200 38548 15252 38554
rect 15200 38490 15252 38496
rect 15396 36786 15424 39578
rect 15580 39098 15608 39986
rect 16684 39982 16712 41074
rect 17960 40928 18012 40934
rect 18156 40905 18184 41074
rect 17960 40870 18012 40876
rect 18142 40896 18198 40905
rect 17408 40384 17460 40390
rect 17408 40326 17460 40332
rect 16672 39976 16724 39982
rect 16672 39918 16724 39924
rect 16120 39908 16172 39914
rect 16120 39850 16172 39856
rect 15776 39740 16084 39760
rect 15776 39738 15782 39740
rect 15838 39738 15862 39740
rect 15918 39738 15942 39740
rect 15998 39738 16022 39740
rect 16078 39738 16084 39740
rect 15838 39686 15840 39738
rect 16020 39686 16022 39738
rect 15776 39684 15782 39686
rect 15838 39684 15862 39686
rect 15918 39684 15942 39686
rect 15998 39684 16022 39686
rect 16078 39684 16084 39686
rect 15776 39664 16084 39684
rect 15752 39568 15804 39574
rect 15752 39510 15804 39516
rect 15660 39432 15712 39438
rect 15660 39374 15712 39380
rect 15568 39092 15620 39098
rect 15568 39034 15620 39040
rect 15672 39030 15700 39374
rect 15660 39024 15712 39030
rect 15660 38966 15712 38972
rect 15764 38962 15792 39510
rect 15936 39296 15988 39302
rect 15936 39238 15988 39244
rect 15948 38962 15976 39238
rect 15752 38956 15804 38962
rect 15752 38898 15804 38904
rect 15936 38956 15988 38962
rect 15936 38898 15988 38904
rect 15776 38652 16084 38672
rect 15776 38650 15782 38652
rect 15838 38650 15862 38652
rect 15918 38650 15942 38652
rect 15998 38650 16022 38652
rect 16078 38650 16084 38652
rect 15838 38598 15840 38650
rect 16020 38598 16022 38650
rect 15776 38596 15782 38598
rect 15838 38596 15862 38598
rect 15918 38596 15942 38598
rect 15998 38596 16022 38598
rect 16078 38596 16084 38598
rect 15776 38576 16084 38596
rect 15776 37564 16084 37584
rect 15776 37562 15782 37564
rect 15838 37562 15862 37564
rect 15918 37562 15942 37564
rect 15998 37562 16022 37564
rect 16078 37562 16084 37564
rect 15838 37510 15840 37562
rect 16020 37510 16022 37562
rect 15776 37508 15782 37510
rect 15838 37508 15862 37510
rect 15918 37508 15942 37510
rect 15998 37508 16022 37510
rect 16078 37508 16084 37510
rect 15776 37488 16084 37508
rect 15384 36780 15436 36786
rect 15384 36722 15436 36728
rect 15568 36780 15620 36786
rect 15568 36722 15620 36728
rect 15384 36576 15436 36582
rect 15384 36518 15436 36524
rect 14924 36168 14976 36174
rect 14924 36110 14976 36116
rect 14740 36032 14792 36038
rect 14740 35974 14792 35980
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 14556 35624 14608 35630
rect 14556 35566 14608 35572
rect 14568 35154 14596 35566
rect 14556 35148 14608 35154
rect 14556 35090 14608 35096
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 14188 34944 14240 34950
rect 14188 34886 14240 34892
rect 14200 34678 14228 34886
rect 14188 34672 14240 34678
rect 14188 34614 14240 34620
rect 14568 34610 14596 35090
rect 14752 35086 14780 35974
rect 15212 35222 15240 35974
rect 15396 35698 15424 36518
rect 15384 35692 15436 35698
rect 15384 35634 15436 35640
rect 15200 35216 15252 35222
rect 15200 35158 15252 35164
rect 14740 35080 14792 35086
rect 14740 35022 14792 35028
rect 14832 35080 14884 35086
rect 14832 35022 14884 35028
rect 14556 34604 14608 34610
rect 14556 34546 14608 34552
rect 14844 34202 14872 35022
rect 15580 34610 15608 36722
rect 15776 36476 16084 36496
rect 15776 36474 15782 36476
rect 15838 36474 15862 36476
rect 15918 36474 15942 36476
rect 15998 36474 16022 36476
rect 16078 36474 16084 36476
rect 15838 36422 15840 36474
rect 16020 36422 16022 36474
rect 15776 36420 15782 36422
rect 15838 36420 15862 36422
rect 15918 36420 15942 36422
rect 15998 36420 16022 36422
rect 16078 36420 16084 36422
rect 15776 36400 16084 36420
rect 16132 36038 16160 39850
rect 17420 36718 17448 40326
rect 17972 39370 18000 40870
rect 18142 40831 18198 40840
rect 17960 39364 18012 39370
rect 17960 39306 18012 39312
rect 16580 36712 16632 36718
rect 16580 36654 16632 36660
rect 17408 36712 17460 36718
rect 17408 36654 17460 36660
rect 16592 36310 16620 36654
rect 16580 36304 16632 36310
rect 16580 36246 16632 36252
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 15660 36032 15712 36038
rect 15660 35974 15712 35980
rect 16120 36032 16172 36038
rect 16172 35992 16344 36020
rect 16120 35974 16172 35980
rect 15672 35494 15700 35974
rect 16316 35494 16344 35992
rect 16500 35834 16528 36110
rect 16764 36032 16816 36038
rect 16764 35974 16816 35980
rect 16488 35828 16540 35834
rect 16488 35770 16540 35776
rect 16776 35630 16804 35974
rect 17420 35698 17448 36654
rect 17408 35692 17460 35698
rect 17408 35634 17460 35640
rect 16764 35624 16816 35630
rect 16764 35566 16816 35572
rect 15660 35488 15712 35494
rect 15660 35430 15712 35436
rect 16304 35488 16356 35494
rect 16304 35430 16356 35436
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 15016 34536 15068 34542
rect 15016 34478 15068 34484
rect 14832 34196 14884 34202
rect 14832 34138 14884 34144
rect 14096 33992 14148 33998
rect 14096 33934 14148 33940
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 14108 33114 14136 33934
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14096 33108 14148 33114
rect 14096 33050 14148 33056
rect 13728 32904 13780 32910
rect 13728 32846 13780 32852
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 13740 32230 13768 32846
rect 13728 32224 13780 32230
rect 13728 32166 13780 32172
rect 13740 30258 13768 32166
rect 14200 31754 14228 32846
rect 14108 31726 14228 31754
rect 14004 30592 14056 30598
rect 14004 30534 14056 30540
rect 14016 30258 14044 30534
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 13728 29844 13780 29850
rect 13728 29786 13780 29792
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13544 28484 13596 28490
rect 13544 28426 13596 28432
rect 13556 27606 13584 28426
rect 13648 28150 13676 29446
rect 13740 28626 13768 29786
rect 13728 28620 13780 28626
rect 13728 28562 13780 28568
rect 13740 28218 13768 28562
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 13544 27600 13596 27606
rect 13544 27542 13596 27548
rect 13832 27402 13860 28426
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 14016 27470 14044 28358
rect 14004 27464 14056 27470
rect 14004 27406 14056 27412
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13452 26852 13504 26858
rect 13452 26794 13504 26800
rect 14108 26382 14136 31726
rect 14384 31346 14412 33458
rect 15028 33454 15056 34478
rect 15672 34066 15700 35430
rect 15776 35388 16084 35408
rect 15776 35386 15782 35388
rect 15838 35386 15862 35388
rect 15918 35386 15942 35388
rect 15998 35386 16022 35388
rect 16078 35386 16084 35388
rect 15838 35334 15840 35386
rect 16020 35334 16022 35386
rect 15776 35332 15782 35334
rect 15838 35332 15862 35334
rect 15918 35332 15942 35334
rect 15998 35332 16022 35334
rect 16078 35332 16084 35334
rect 15776 35312 16084 35332
rect 16776 35290 16804 35566
rect 16764 35284 16816 35290
rect 16764 35226 16816 35232
rect 16672 35012 16724 35018
rect 16672 34954 16724 34960
rect 16304 34944 16356 34950
rect 16304 34886 16356 34892
rect 15776 34300 16084 34320
rect 15776 34298 15782 34300
rect 15838 34298 15862 34300
rect 15918 34298 15942 34300
rect 15998 34298 16022 34300
rect 16078 34298 16084 34300
rect 15838 34246 15840 34298
rect 16020 34246 16022 34298
rect 15776 34244 15782 34246
rect 15838 34244 15862 34246
rect 15918 34244 15942 34246
rect 15998 34244 16022 34246
rect 16078 34244 16084 34246
rect 15776 34224 16084 34244
rect 15660 34060 15712 34066
rect 15660 34002 15712 34008
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 15016 33448 15068 33454
rect 15016 33390 15068 33396
rect 15028 32910 15056 33390
rect 15396 32978 15424 33866
rect 15776 33212 16084 33232
rect 15776 33210 15782 33212
rect 15838 33210 15862 33212
rect 15918 33210 15942 33212
rect 15998 33210 16022 33212
rect 16078 33210 16084 33212
rect 15838 33158 15840 33210
rect 16020 33158 16022 33210
rect 15776 33156 15782 33158
rect 15838 33156 15862 33158
rect 15918 33156 15942 33158
rect 15998 33156 16022 33158
rect 16078 33156 16084 33158
rect 15776 33136 16084 33156
rect 15384 32972 15436 32978
rect 15384 32914 15436 32920
rect 15016 32904 15068 32910
rect 15016 32846 15068 32852
rect 14188 31340 14240 31346
rect 14188 31282 14240 31288
rect 14372 31340 14424 31346
rect 14372 31282 14424 31288
rect 14200 29714 14228 31282
rect 14280 31272 14332 31278
rect 14280 31214 14332 31220
rect 14292 30598 14320 31214
rect 14280 30592 14332 30598
rect 14280 30534 14332 30540
rect 14188 29708 14240 29714
rect 14188 29650 14240 29656
rect 14292 29646 14320 30534
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14476 29782 14504 30194
rect 14464 29776 14516 29782
rect 14464 29718 14516 29724
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14292 28694 14320 29582
rect 14384 29306 14412 29582
rect 14556 29572 14608 29578
rect 14556 29514 14608 29520
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14280 28688 14332 28694
rect 14280 28630 14332 28636
rect 14384 28558 14412 29242
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14568 28490 14596 29514
rect 14556 28484 14608 28490
rect 14556 28426 14608 28432
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14292 27674 14320 28018
rect 14280 27668 14332 27674
rect 14280 27610 14332 27616
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 12811 26140 13119 26160
rect 12811 26138 12817 26140
rect 12873 26138 12897 26140
rect 12953 26138 12977 26140
rect 13033 26138 13057 26140
rect 13113 26138 13119 26140
rect 12873 26086 12875 26138
rect 13055 26086 13057 26138
rect 12811 26084 12817 26086
rect 12873 26084 12897 26086
rect 12953 26084 12977 26086
rect 13033 26084 13057 26086
rect 13113 26084 13119 26086
rect 12811 26064 13119 26084
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12820 25498 12848 25842
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12544 24954 12572 25230
rect 12811 25052 13119 25072
rect 12811 25050 12817 25052
rect 12873 25050 12897 25052
rect 12953 25050 12977 25052
rect 13033 25050 13057 25052
rect 13113 25050 13119 25052
rect 12873 24998 12875 25050
rect 13055 24998 13057 25050
rect 12811 24996 12817 24998
rect 12873 24996 12897 24998
rect 12953 24996 12977 24998
rect 13033 24996 13057 24998
rect 13113 24996 13119 24998
rect 12811 24976 13119 24996
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12268 23798 12296 24550
rect 14108 24206 14136 26318
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14476 24954 14504 25230
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14464 24948 14516 24954
rect 14464 24890 14516 24896
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 12811 23964 13119 23984
rect 12811 23962 12817 23964
rect 12873 23962 12897 23964
rect 12953 23962 12977 23964
rect 13033 23962 13057 23964
rect 13113 23962 13119 23964
rect 12873 23910 12875 23962
rect 13055 23910 13057 23962
rect 12811 23908 12817 23910
rect 12873 23908 12897 23910
rect 12953 23908 12977 23910
rect 13033 23908 13057 23910
rect 13113 23908 13119 23910
rect 12811 23888 13119 23908
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12268 22574 12296 23734
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 13280 23118 13308 23462
rect 13648 23254 13676 23598
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13636 23248 13688 23254
rect 13636 23190 13688 23196
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12084 22066 12204 22094
rect 12176 20330 12204 22066
rect 12544 21690 12572 22578
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12084 18222 12112 18702
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12084 16250 12112 18158
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 12084 14822 12112 15370
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12084 14346 12112 14758
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12176 12306 12204 20266
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12452 18290 12480 18702
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12268 17746 12296 18022
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12268 17202 12296 17682
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12360 17270 12388 17546
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12268 16726 12296 17002
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12360 16182 12388 16730
rect 12452 16454 12480 18226
rect 12544 17678 12572 18838
rect 12636 17882 12664 22918
rect 12811 22876 13119 22896
rect 12811 22874 12817 22876
rect 12873 22874 12897 22876
rect 12953 22874 12977 22876
rect 13033 22874 13057 22876
rect 13113 22874 13119 22876
rect 12873 22822 12875 22874
rect 13055 22822 13057 22874
rect 12811 22820 12817 22822
rect 12873 22820 12897 22822
rect 12953 22820 12977 22822
rect 13033 22820 13057 22822
rect 13113 22820 13119 22822
rect 12811 22800 13119 22820
rect 13188 22778 13216 23054
rect 13176 22772 13228 22778
rect 13176 22714 13228 22720
rect 13188 22094 13216 22714
rect 13280 22234 13308 23054
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 13360 22160 13412 22166
rect 13360 22102 13412 22108
rect 13188 22066 13308 22094
rect 13280 22030 13308 22066
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 12811 21788 13119 21808
rect 12811 21786 12817 21788
rect 12873 21786 12897 21788
rect 12953 21786 12977 21788
rect 13033 21786 13057 21788
rect 13113 21786 13119 21788
rect 12873 21734 12875 21786
rect 13055 21734 13057 21786
rect 12811 21732 12817 21734
rect 12873 21732 12897 21734
rect 12953 21732 12977 21734
rect 13033 21732 13057 21734
rect 13113 21732 13119 21734
rect 12811 21712 13119 21732
rect 13372 20942 13400 22102
rect 13464 22098 13492 23122
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22098 13584 22918
rect 13648 22506 13676 23190
rect 13832 23118 13860 23462
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13636 22500 13688 22506
rect 13636 22442 13688 22448
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13544 22092 13596 22098
rect 14476 22094 14504 24142
rect 14556 23248 14608 23254
rect 14556 23190 14608 23196
rect 14568 22574 14596 23190
rect 14660 23050 14688 24686
rect 14844 23730 14872 25094
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 13544 22034 13596 22040
rect 14384 22066 14504 22094
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13464 21554 13492 21830
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 12728 20466 12756 20878
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 12811 20700 13119 20720
rect 12811 20698 12817 20700
rect 12873 20698 12897 20700
rect 12953 20698 12977 20700
rect 13033 20698 13057 20700
rect 13113 20698 13119 20700
rect 12873 20646 12875 20698
rect 13055 20646 13057 20698
rect 12811 20644 12817 20646
rect 12873 20644 12897 20646
rect 12953 20644 12977 20646
rect 13033 20644 13057 20646
rect 13113 20644 13119 20646
rect 12811 20624 13119 20644
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12728 19786 12756 20402
rect 12716 19780 12768 19786
rect 12716 19722 12768 19728
rect 12728 19378 12756 19722
rect 12811 19612 13119 19632
rect 12811 19610 12817 19612
rect 12873 19610 12897 19612
rect 12953 19610 12977 19612
rect 13033 19610 13057 19612
rect 13113 19610 13119 19612
rect 12873 19558 12875 19610
rect 13055 19558 13057 19610
rect 12811 19556 12817 19558
rect 12873 19556 12897 19558
rect 12953 19556 12977 19558
rect 13033 19556 13057 19558
rect 13113 19556 13119 19558
rect 12811 19536 13119 19556
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12728 17814 12756 19314
rect 13188 19174 13216 20742
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13188 18834 13216 19110
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13372 18766 13400 19246
rect 13360 18760 13412 18766
rect 13412 18720 13492 18748
rect 13360 18702 13412 18708
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 12811 18524 13119 18544
rect 12811 18522 12817 18524
rect 12873 18522 12897 18524
rect 12953 18522 12977 18524
rect 13033 18522 13057 18524
rect 13113 18522 13119 18524
rect 12873 18470 12875 18522
rect 13055 18470 13057 18522
rect 12811 18468 12817 18470
rect 12873 18468 12897 18470
rect 12953 18468 12977 18470
rect 13033 18468 13057 18470
rect 13113 18468 13119 18470
rect 12811 18448 13119 18468
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 13372 17678 13400 18566
rect 12532 17672 12584 17678
rect 12808 17672 12860 17678
rect 12584 17632 12664 17660
rect 12532 17614 12584 17620
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12544 15502 12572 17478
rect 12636 16998 12664 17632
rect 12728 17632 12808 17660
rect 12728 17066 12756 17632
rect 12808 17614 12860 17620
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 12811 17436 13119 17456
rect 12811 17434 12817 17436
rect 12873 17434 12897 17436
rect 12953 17434 12977 17436
rect 13033 17434 13057 17436
rect 13113 17434 13119 17436
rect 12873 17382 12875 17434
rect 13055 17382 13057 17434
rect 12811 17380 12817 17382
rect 12873 17380 12897 17382
rect 12953 17380 12977 17382
rect 13033 17380 13057 17382
rect 13113 17380 13119 17382
rect 12811 17360 13119 17380
rect 13464 17202 13492 18720
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12728 12442 12756 17002
rect 13280 16726 13308 17070
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 12811 16348 13119 16368
rect 12811 16346 12817 16348
rect 12873 16346 12897 16348
rect 12953 16346 12977 16348
rect 13033 16346 13057 16348
rect 13113 16346 13119 16348
rect 12873 16294 12875 16346
rect 13055 16294 13057 16346
rect 12811 16292 12817 16294
rect 12873 16292 12897 16294
rect 12953 16292 12977 16294
rect 13033 16292 13057 16294
rect 13113 16292 13119 16294
rect 12811 16272 13119 16292
rect 12811 15260 13119 15280
rect 12811 15258 12817 15260
rect 12873 15258 12897 15260
rect 12953 15258 12977 15260
rect 13033 15258 13057 15260
rect 13113 15258 13119 15260
rect 12873 15206 12875 15258
rect 13055 15206 13057 15258
rect 12811 15204 12817 15206
rect 12873 15204 12897 15206
rect 12953 15204 12977 15206
rect 13033 15204 13057 15206
rect 13113 15204 13119 15206
rect 12811 15184 13119 15204
rect 12811 14172 13119 14192
rect 12811 14170 12817 14172
rect 12873 14170 12897 14172
rect 12953 14170 12977 14172
rect 13033 14170 13057 14172
rect 13113 14170 13119 14172
rect 12873 14118 12875 14170
rect 13055 14118 13057 14170
rect 12811 14116 12817 14118
rect 12873 14116 12897 14118
rect 12953 14116 12977 14118
rect 13033 14116 13057 14118
rect 13113 14116 13119 14118
rect 12811 14096 13119 14116
rect 12811 13084 13119 13104
rect 12811 13082 12817 13084
rect 12873 13082 12897 13084
rect 12953 13082 12977 13084
rect 13033 13082 13057 13084
rect 13113 13082 13119 13084
rect 12873 13030 12875 13082
rect 13055 13030 13057 13082
rect 12811 13028 12817 13030
rect 12873 13028 12897 13030
rect 12953 13028 12977 13030
rect 13033 13028 13057 13030
rect 13113 13028 13119 13030
rect 12811 13008 13119 13028
rect 13280 12986 13308 16662
rect 13464 16658 13492 17002
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13556 14550 13584 21898
rect 14384 19310 14412 22066
rect 14568 22030 14596 22510
rect 14660 22506 14688 22986
rect 15028 22642 15056 32846
rect 15776 32124 16084 32144
rect 15776 32122 15782 32124
rect 15838 32122 15862 32124
rect 15918 32122 15942 32124
rect 15998 32122 16022 32124
rect 16078 32122 16084 32124
rect 15838 32070 15840 32122
rect 16020 32070 16022 32122
rect 15776 32068 15782 32070
rect 15838 32068 15862 32070
rect 15918 32068 15942 32070
rect 15998 32068 16022 32070
rect 16078 32068 16084 32070
rect 15776 32048 16084 32068
rect 16210 32056 16266 32065
rect 16132 32014 16210 32042
rect 15776 31036 16084 31056
rect 15776 31034 15782 31036
rect 15838 31034 15862 31036
rect 15918 31034 15942 31036
rect 15998 31034 16022 31036
rect 16078 31034 16084 31036
rect 15838 30982 15840 31034
rect 16020 30982 16022 31034
rect 15776 30980 15782 30982
rect 15838 30980 15862 30982
rect 15918 30980 15942 30982
rect 15998 30980 16022 30982
rect 16078 30980 16084 30982
rect 15776 30960 16084 30980
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15488 30326 15516 30670
rect 15752 30660 15804 30666
rect 15752 30602 15804 30608
rect 15764 30394 15792 30602
rect 15752 30388 15804 30394
rect 15752 30330 15804 30336
rect 15476 30320 15528 30326
rect 15476 30262 15528 30268
rect 15108 30048 15160 30054
rect 15108 29990 15160 29996
rect 15120 29646 15148 29990
rect 15488 29714 15516 30262
rect 15776 29948 16084 29968
rect 15776 29946 15782 29948
rect 15838 29946 15862 29948
rect 15918 29946 15942 29948
rect 15998 29946 16022 29948
rect 16078 29946 16084 29948
rect 15838 29894 15840 29946
rect 16020 29894 16022 29946
rect 15776 29892 15782 29894
rect 15838 29892 15862 29894
rect 15918 29892 15942 29894
rect 15998 29892 16022 29894
rect 16078 29892 16084 29894
rect 15776 29872 16084 29892
rect 15476 29708 15528 29714
rect 15476 29650 15528 29656
rect 15108 29640 15160 29646
rect 15108 29582 15160 29588
rect 15488 29170 15516 29650
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 15856 29170 15884 29446
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 15488 28626 15516 29106
rect 15776 28860 16084 28880
rect 15776 28858 15782 28860
rect 15838 28858 15862 28860
rect 15918 28858 15942 28860
rect 15998 28858 16022 28860
rect 16078 28858 16084 28860
rect 15838 28806 15840 28858
rect 16020 28806 16022 28858
rect 15776 28804 15782 28806
rect 15838 28804 15862 28806
rect 15918 28804 15942 28806
rect 15998 28804 16022 28806
rect 16078 28804 16084 28806
rect 15776 28784 16084 28804
rect 15476 28620 15528 28626
rect 15476 28562 15528 28568
rect 15488 28082 15516 28562
rect 15476 28076 15528 28082
rect 15476 28018 15528 28024
rect 15776 27772 16084 27792
rect 15776 27770 15782 27772
rect 15838 27770 15862 27772
rect 15918 27770 15942 27772
rect 15998 27770 16022 27772
rect 16078 27770 16084 27772
rect 15838 27718 15840 27770
rect 16020 27718 16022 27770
rect 15776 27716 15782 27718
rect 15838 27716 15862 27718
rect 15918 27716 15942 27718
rect 15998 27716 16022 27718
rect 16078 27716 16084 27718
rect 15776 27696 16084 27716
rect 15776 26684 16084 26704
rect 15776 26682 15782 26684
rect 15838 26682 15862 26684
rect 15918 26682 15942 26684
rect 15998 26682 16022 26684
rect 16078 26682 16084 26684
rect 15838 26630 15840 26682
rect 16020 26630 16022 26682
rect 15776 26628 15782 26630
rect 15838 26628 15862 26630
rect 15918 26628 15942 26630
rect 15998 26628 16022 26630
rect 16078 26628 16084 26630
rect 15776 26608 16084 26628
rect 15476 25900 15528 25906
rect 15476 25842 15528 25848
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15304 24818 15332 25094
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15108 24608 15160 24614
rect 15160 24568 15240 24596
rect 15108 24550 15160 24556
rect 15212 24206 15240 24568
rect 15488 24410 15516 25842
rect 15568 25696 15620 25702
rect 15568 25638 15620 25644
rect 15580 25294 15608 25638
rect 15776 25596 16084 25616
rect 15776 25594 15782 25596
rect 15838 25594 15862 25596
rect 15918 25594 15942 25596
rect 15998 25594 16022 25596
rect 16078 25594 16084 25596
rect 15838 25542 15840 25594
rect 16020 25542 16022 25594
rect 15776 25540 15782 25542
rect 15838 25540 15862 25542
rect 15918 25540 15942 25542
rect 15998 25540 16022 25542
rect 16078 25540 16084 25542
rect 15776 25520 16084 25540
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15212 23798 15240 24142
rect 15580 24138 15608 25230
rect 15776 24508 16084 24528
rect 15776 24506 15782 24508
rect 15838 24506 15862 24508
rect 15918 24506 15942 24508
rect 15998 24506 16022 24508
rect 16078 24506 16084 24508
rect 15838 24454 15840 24506
rect 16020 24454 16022 24506
rect 15776 24452 15782 24454
rect 15838 24452 15862 24454
rect 15918 24452 15942 24454
rect 15998 24452 16022 24454
rect 16078 24452 16084 24454
rect 15776 24432 16084 24452
rect 15568 24132 15620 24138
rect 15568 24074 15620 24080
rect 16132 24070 16160 32014
rect 16210 31991 16266 32000
rect 16316 25430 16344 34886
rect 16684 34746 16712 34954
rect 16672 34740 16724 34746
rect 16672 34682 16724 34688
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 16868 34202 16896 34546
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16764 32972 16816 32978
rect 16764 32914 16816 32920
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16592 30190 16620 30534
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16592 25906 16620 30126
rect 16684 29578 16712 31078
rect 16776 30258 16804 32914
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16868 30394 16896 31282
rect 17500 30660 17552 30666
rect 17500 30602 17552 30608
rect 17512 30394 17540 30602
rect 16856 30388 16908 30394
rect 16856 30330 16908 30336
rect 17500 30388 17552 30394
rect 17500 30330 17552 30336
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 17684 30252 17736 30258
rect 17684 30194 17736 30200
rect 16672 29572 16724 29578
rect 16672 29514 16724 29520
rect 16960 29170 16988 30194
rect 17592 29504 17644 29510
rect 17592 29446 17644 29452
rect 16764 29164 16816 29170
rect 16764 29106 16816 29112
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 16776 28762 16804 29106
rect 16764 28756 16816 28762
rect 16764 28698 16816 28704
rect 16672 28484 16724 28490
rect 16672 28426 16724 28432
rect 16684 28218 16712 28426
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 16776 27146 16804 28698
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16684 27118 16804 27146
rect 16868 27130 16896 28018
rect 16856 27124 16908 27130
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16304 25424 16356 25430
rect 16304 25366 16356 25372
rect 16316 25226 16344 25366
rect 16592 25362 16620 25842
rect 16684 25498 16712 27118
rect 16856 27066 16908 27072
rect 16960 26994 16988 29106
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16776 25838 16804 26930
rect 16764 25832 16816 25838
rect 16764 25774 16816 25780
rect 16672 25492 16724 25498
rect 16672 25434 16724 25440
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 16684 24818 16712 25230
rect 16776 25226 16804 25774
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16776 24410 16804 25162
rect 16868 24818 16896 25434
rect 16960 24954 16988 26930
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 16948 24948 17000 24954
rect 16948 24890 17000 24896
rect 17052 24818 17080 25638
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17144 24410 17172 25094
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 16764 24404 16816 24410
rect 16764 24346 16816 24352
rect 17132 24404 17184 24410
rect 17132 24346 17184 24352
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16120 24064 16172 24070
rect 16120 24006 16172 24012
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 15776 23420 16084 23440
rect 15776 23418 15782 23420
rect 15838 23418 15862 23420
rect 15918 23418 15942 23420
rect 15998 23418 16022 23420
rect 16078 23418 16084 23420
rect 15838 23366 15840 23418
rect 16020 23366 16022 23418
rect 15776 23364 15782 23366
rect 15838 23364 15862 23366
rect 15918 23364 15942 23366
rect 15998 23364 16022 23366
rect 16078 23364 16084 23366
rect 15776 23344 16084 23364
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 16040 22642 16068 23054
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 14648 22500 14700 22506
rect 14648 22442 14700 22448
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 14108 17678 14136 18294
rect 14568 18086 14596 21966
rect 15028 19990 15056 22578
rect 15672 22098 15700 22578
rect 15776 22332 16084 22352
rect 15776 22330 15782 22332
rect 15838 22330 15862 22332
rect 15918 22330 15942 22332
rect 15998 22330 16022 22332
rect 16078 22330 16084 22332
rect 15838 22278 15840 22330
rect 16020 22278 16022 22330
rect 15776 22276 15782 22278
rect 15838 22276 15862 22278
rect 15918 22276 15942 22278
rect 15998 22276 16022 22278
rect 16078 22276 16084 22278
rect 15776 22256 16084 22276
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15016 19984 15068 19990
rect 15016 19926 15068 19932
rect 15028 19378 15056 19926
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15120 19446 15148 19790
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 15120 18970 15148 19382
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14936 18290 14964 18702
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 16794 14136 17614
rect 14660 17338 14688 18226
rect 15120 17882 15148 18906
rect 15212 18358 15240 19450
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 15304 18290 15332 20470
rect 15672 19854 15700 22034
rect 15776 21244 16084 21264
rect 15776 21242 15782 21244
rect 15838 21242 15862 21244
rect 15918 21242 15942 21244
rect 15998 21242 16022 21244
rect 16078 21242 16084 21244
rect 15838 21190 15840 21242
rect 16020 21190 16022 21242
rect 15776 21188 15782 21190
rect 15838 21188 15862 21190
rect 15918 21188 15942 21190
rect 15998 21188 16022 21190
rect 16078 21188 16084 21190
rect 15776 21168 16084 21188
rect 16132 21146 16160 23666
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16224 23225 16252 23462
rect 16210 23216 16266 23225
rect 16592 23186 16620 24074
rect 17420 24070 17448 24686
rect 17604 24614 17632 29446
rect 17696 29306 17724 30194
rect 17684 29300 17736 29306
rect 17684 29242 17736 29248
rect 17960 25764 18012 25770
rect 17960 25706 18012 25712
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17604 24138 17632 24550
rect 17972 24290 18000 25706
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17880 24274 18000 24290
rect 17868 24268 18000 24274
rect 17920 24262 18000 24268
rect 17868 24210 17920 24216
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17420 23866 17448 24006
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 16776 23186 16804 23666
rect 16210 23151 16266 23160
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16776 22642 16804 23122
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 16948 22976 17000 22982
rect 16948 22918 17000 22924
rect 16960 22794 16988 22918
rect 16960 22766 17080 22794
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 16960 22386 16988 22578
rect 16776 22358 16988 22386
rect 16776 21894 16804 22358
rect 17052 22094 17080 22766
rect 16960 22066 17080 22094
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 16960 21554 16988 22066
rect 17144 21690 17172 22986
rect 17604 21690 17632 23666
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 17788 21554 17816 21830
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15776 20156 16084 20176
rect 15776 20154 15782 20156
rect 15838 20154 15862 20156
rect 15918 20154 15942 20156
rect 15998 20154 16022 20156
rect 16078 20154 16084 20156
rect 15838 20102 15840 20154
rect 16020 20102 16022 20154
rect 15776 20100 15782 20102
rect 15838 20100 15862 20102
rect 15918 20100 15942 20102
rect 15998 20100 16022 20102
rect 16078 20100 16084 20102
rect 15776 20080 16084 20100
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16684 19378 16712 19654
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 15384 19236 15436 19242
rect 15384 19178 15436 19184
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14844 17202 14872 17546
rect 15212 17202 15240 18022
rect 15396 17814 15424 19178
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 15776 19068 16084 19088
rect 15776 19066 15782 19068
rect 15838 19066 15862 19068
rect 15918 19066 15942 19068
rect 15998 19066 16022 19068
rect 16078 19066 16084 19068
rect 15838 19014 15840 19066
rect 16020 19014 16022 19066
rect 15776 19012 15782 19014
rect 15838 19012 15862 19014
rect 15918 19012 15942 19014
rect 15998 19012 16022 19014
rect 16078 19012 16084 19014
rect 15776 18992 16084 19012
rect 16132 18970 16160 19110
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15384 17808 15436 17814
rect 15384 17750 15436 17756
rect 15488 17338 15516 18634
rect 15776 17980 16084 18000
rect 15776 17978 15782 17980
rect 15838 17978 15862 17980
rect 15918 17978 15942 17980
rect 15998 17978 16022 17980
rect 16078 17978 16084 17980
rect 15838 17926 15840 17978
rect 16020 17926 16022 17978
rect 15776 17924 15782 17926
rect 15838 17924 15862 17926
rect 15918 17924 15942 17926
rect 15998 17924 16022 17926
rect 16078 17924 16084 17926
rect 15776 17904 16084 17924
rect 16132 17678 16160 18906
rect 16224 18290 16252 19246
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16224 17746 16252 18226
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16120 17672 16172 17678
rect 16040 17632 16120 17660
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15948 17270 15976 17478
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 16040 17134 16068 17632
rect 16120 17614 16172 17620
rect 16316 17610 16344 18158
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 15028 16590 15056 16934
rect 15776 16892 16084 16912
rect 15776 16890 15782 16892
rect 15838 16890 15862 16892
rect 15918 16890 15942 16892
rect 15998 16890 16022 16892
rect 16078 16890 16084 16892
rect 15838 16838 15840 16890
rect 16020 16838 16022 16890
rect 15776 16836 15782 16838
rect 15838 16836 15862 16838
rect 15918 16836 15942 16838
rect 15998 16836 16022 16838
rect 16078 16836 16084 16838
rect 15776 16816 16084 16836
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 14384 15434 14412 16458
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14844 16046 14872 16390
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 14384 14006 14412 15370
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13372 12646 13400 13806
rect 13832 13326 13860 13874
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12084 10742 12112 11154
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11992 8634 12020 9998
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11808 7342 11836 8434
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11532 3738 11560 5170
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4622 11744 4966
rect 11808 4826 11836 7278
rect 11900 5914 11928 7346
rect 11992 7206 12020 8434
rect 12084 7886 12112 10678
rect 12176 10130 12204 12242
rect 13372 12102 13400 12582
rect 13464 12170 13492 13194
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 12811 11996 13119 12016
rect 12811 11994 12817 11996
rect 12873 11994 12897 11996
rect 12953 11994 12977 11996
rect 13033 11994 13057 11996
rect 13113 11994 13119 11996
rect 12873 11942 12875 11994
rect 13055 11942 13057 11994
rect 12811 11940 12817 11942
rect 12873 11940 12897 11942
rect 12953 11940 12977 11942
rect 13033 11940 13057 11942
rect 13113 11940 13119 11942
rect 12811 11920 13119 11940
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12544 9722 12572 10542
rect 12728 10266 12756 11698
rect 13188 11354 13216 12038
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13372 11082 13400 12038
rect 13464 11558 13492 12106
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11150 13492 11494
rect 13556 11218 13584 13262
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13740 12442 13768 12786
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 12811 10908 13119 10928
rect 12811 10906 12817 10908
rect 12873 10906 12897 10908
rect 12953 10906 12977 10908
rect 13033 10906 13057 10908
rect 13113 10906 13119 10908
rect 12873 10854 12875 10906
rect 13055 10854 13057 10906
rect 12811 10852 12817 10854
rect 12873 10852 12897 10854
rect 12953 10852 12977 10854
rect 13033 10852 13057 10854
rect 13113 10852 13119 10854
rect 12811 10832 13119 10852
rect 13556 10674 13584 11154
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12912 10062 12940 10406
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12811 9820 13119 9840
rect 12811 9818 12817 9820
rect 12873 9818 12897 9820
rect 12953 9818 12977 9820
rect 13033 9818 13057 9820
rect 13113 9818 13119 9820
rect 12873 9766 12875 9818
rect 13055 9766 13057 9818
rect 12811 9764 12817 9766
rect 12873 9764 12897 9766
rect 12953 9764 12977 9766
rect 13033 9764 13057 9766
rect 13113 9764 13119 9766
rect 12811 9744 13119 9764
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6798 12480 7142
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 6458 12480 6598
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 12176 5642 12204 6258
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12268 5710 12296 6122
rect 12452 5778 12480 6394
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12176 5370 12204 5578
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12268 5250 12296 5646
rect 12176 5222 12296 5250
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 12176 3942 12204 5222
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 12544 3670 12572 9658
rect 12811 8732 13119 8752
rect 12811 8730 12817 8732
rect 12873 8730 12897 8732
rect 12953 8730 12977 8732
rect 13033 8730 13057 8732
rect 13113 8730 13119 8732
rect 12873 8678 12875 8730
rect 13055 8678 13057 8730
rect 12811 8676 12817 8678
rect 12873 8676 12897 8678
rect 12953 8676 12977 8678
rect 13033 8676 13057 8678
rect 13113 8676 13119 8678
rect 12811 8656 13119 8676
rect 13188 8498 13216 10610
rect 13740 10606 13768 11290
rect 13832 10674 13860 13126
rect 14108 12238 14136 13126
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14200 12306 14228 12378
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 12811 7644 13119 7664
rect 12811 7642 12817 7644
rect 12873 7642 12897 7644
rect 12953 7642 12977 7644
rect 13033 7642 13057 7644
rect 13113 7642 13119 7644
rect 12873 7590 12875 7642
rect 13055 7590 13057 7642
rect 12811 7588 12817 7590
rect 12873 7588 12897 7590
rect 12953 7588 12977 7590
rect 13033 7588 13057 7590
rect 13113 7588 13119 7590
rect 12811 7568 13119 7588
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12636 6458 12664 7346
rect 12811 6556 13119 6576
rect 12811 6554 12817 6556
rect 12873 6554 12897 6556
rect 12953 6554 12977 6556
rect 13033 6554 13057 6556
rect 13113 6554 13119 6556
rect 12873 6502 12875 6554
rect 13055 6502 13057 6554
rect 12811 6500 12817 6502
rect 12873 6500 12897 6502
rect 12953 6500 12977 6502
rect 13033 6500 13057 6502
rect 13113 6500 13119 6502
rect 12811 6480 13119 6500
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 13372 6322 13400 7686
rect 13556 7478 13584 7686
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 12636 5914 12664 6258
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12636 4826 12664 5850
rect 13372 5710 13400 6258
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 12811 5468 13119 5488
rect 12811 5466 12817 5468
rect 12873 5466 12897 5468
rect 12953 5466 12977 5468
rect 13033 5466 13057 5468
rect 13113 5466 13119 5468
rect 12873 5414 12875 5466
rect 13055 5414 13057 5466
rect 12811 5412 12817 5414
rect 12873 5412 12897 5414
rect 12953 5412 12977 5414
rect 13033 5412 13057 5414
rect 13113 5412 13119 5414
rect 12811 5392 13119 5412
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 13372 4622 13400 5510
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13464 4826 13492 5170
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 12811 4380 13119 4400
rect 12811 4378 12817 4380
rect 12873 4378 12897 4380
rect 12953 4378 12977 4380
rect 13033 4378 13057 4380
rect 13113 4378 13119 4380
rect 12873 4326 12875 4378
rect 13055 4326 13057 4378
rect 12811 4324 12817 4326
rect 12873 4324 12897 4326
rect 12953 4324 12977 4326
rect 13033 4324 13057 4326
rect 13113 4324 13119 4326
rect 12811 4304 13119 4324
rect 13280 4214 13308 4422
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13740 4010 13768 10542
rect 14016 7342 14044 11630
rect 14108 11218 14136 12174
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14108 7886 14136 8230
rect 14200 8090 14228 11698
rect 14292 10810 14320 12786
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14476 10674 14504 13806
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14752 13326 14780 13738
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14568 11898 14596 12106
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14568 11354 14596 11698
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14660 10810 14688 13194
rect 14752 12850 14780 13262
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14752 12374 14780 12786
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14752 11694 14780 12310
rect 14844 12238 14872 15982
rect 15776 15804 16084 15824
rect 15776 15802 15782 15804
rect 15838 15802 15862 15804
rect 15918 15802 15942 15804
rect 15998 15802 16022 15804
rect 16078 15802 16084 15804
rect 15838 15750 15840 15802
rect 16020 15750 16022 15802
rect 15776 15748 15782 15750
rect 15838 15748 15862 15750
rect 15918 15748 15942 15750
rect 15998 15748 16022 15750
rect 16078 15748 16084 15750
rect 15776 15728 16084 15748
rect 15776 14716 16084 14736
rect 15776 14714 15782 14716
rect 15838 14714 15862 14716
rect 15918 14714 15942 14716
rect 15998 14714 16022 14716
rect 16078 14714 16084 14716
rect 15838 14662 15840 14714
rect 16020 14662 16022 14714
rect 15776 14660 15782 14662
rect 15838 14660 15862 14662
rect 15918 14660 15942 14662
rect 15998 14660 16022 14662
rect 16078 14660 16084 14662
rect 15776 14640 16084 14660
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14752 11150 14780 11630
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14660 7818 14688 8366
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 6798 14044 7278
rect 14660 6914 14688 7754
rect 14752 6934 14780 7822
rect 14568 6886 14688 6914
rect 14740 6928 14792 6934
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14016 5234 14044 6734
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14384 5710 14412 6666
rect 14568 6662 14596 6886
rect 14740 6870 14792 6876
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6458 14596 6598
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14752 5778 14780 6870
rect 14844 6866 14872 12038
rect 15028 11830 15056 14214
rect 15580 14074 15608 14350
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15672 13258 15700 13806
rect 15776 13628 16084 13648
rect 15776 13626 15782 13628
rect 15838 13626 15862 13628
rect 15918 13626 15942 13628
rect 15998 13626 16022 13628
rect 16078 13626 16084 13628
rect 15838 13574 15840 13626
rect 16020 13574 16022 13626
rect 15776 13572 15782 13574
rect 15838 13572 15862 13574
rect 15918 13572 15942 13574
rect 15998 13572 16022 13574
rect 16078 13572 16084 13574
rect 15776 13552 16084 13572
rect 16132 13530 16160 17478
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 13530 16344 16390
rect 16408 13938 16436 17682
rect 16684 17338 16712 18022
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16776 17202 16804 18702
rect 16868 18698 16896 19110
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 16776 16794 16804 17138
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 17328 16250 17356 17138
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 15672 11354 15700 13194
rect 16224 13190 16252 13330
rect 16316 13326 16344 13466
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 15776 12540 16084 12560
rect 15776 12538 15782 12540
rect 15838 12538 15862 12540
rect 15918 12538 15942 12540
rect 15998 12538 16022 12540
rect 16078 12538 16084 12540
rect 15838 12486 15840 12538
rect 16020 12486 16022 12538
rect 15776 12484 15782 12486
rect 15838 12484 15862 12486
rect 15918 12484 15942 12486
rect 15998 12484 16022 12486
rect 16078 12484 16084 12486
rect 15776 12464 16084 12484
rect 16224 11898 16252 13126
rect 16316 12782 16344 13262
rect 16408 12850 16436 13874
rect 17420 13530 17448 18090
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 16590 17632 17478
rect 17972 17338 18000 24262
rect 18064 24138 18092 24754
rect 18156 24206 18184 24754
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 18064 22982 18092 24074
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 18064 21962 18092 22918
rect 18156 22438 18184 24142
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 18156 22098 18184 22374
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18052 21956 18104 21962
rect 18052 21898 18104 21904
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17512 15162 17540 16050
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16684 12782 16712 13262
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16684 12442 16712 12718
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 17420 12238 17448 12582
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17512 12170 17540 12582
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 15776 11452 16084 11472
rect 15776 11450 15782 11452
rect 15838 11450 15862 11452
rect 15918 11450 15942 11452
rect 15998 11450 16022 11452
rect 16078 11450 16084 11452
rect 15838 11398 15840 11450
rect 16020 11398 16022 11450
rect 15776 11396 15782 11398
rect 15838 11396 15862 11398
rect 15918 11396 15942 11398
rect 15998 11396 16022 11398
rect 16078 11396 16084 11398
rect 15776 11376 16084 11396
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14936 6882 14964 8026
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 15396 7206 15424 7890
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 14936 6866 15056 6882
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14936 6860 15068 6866
rect 14936 6854 15016 6860
rect 14936 6730 14964 6854
rect 15016 6802 15068 6808
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 15120 6458 15148 6734
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14016 4146 14044 5170
rect 14292 4622 14320 5510
rect 14752 5370 14780 5714
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14752 4826 14780 5170
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14936 4622 14964 5510
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15120 4146 15148 6394
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15396 4214 15424 4422
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15488 4146 15516 11222
rect 17236 11082 17264 12038
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 15776 10364 16084 10384
rect 15776 10362 15782 10364
rect 15838 10362 15862 10364
rect 15918 10362 15942 10364
rect 15998 10362 16022 10364
rect 16078 10362 16084 10364
rect 15838 10310 15840 10362
rect 16020 10310 16022 10362
rect 15776 10308 15782 10310
rect 15838 10308 15862 10310
rect 15918 10308 15942 10310
rect 15998 10308 16022 10310
rect 16078 10308 16084 10310
rect 15776 10288 16084 10308
rect 17880 9722 17908 14894
rect 17972 14618 18000 14962
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18144 14408 18196 14414
rect 18142 14376 18144 14385
rect 18196 14376 18198 14385
rect 18142 14311 18198 14320
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 15776 9276 16084 9296
rect 15776 9274 15782 9276
rect 15838 9274 15862 9276
rect 15918 9274 15942 9276
rect 15998 9274 16022 9276
rect 16078 9274 16084 9276
rect 15838 9222 15840 9274
rect 16020 9222 16022 9274
rect 15776 9220 15782 9222
rect 15838 9220 15862 9222
rect 15918 9220 15942 9222
rect 15998 9220 16022 9222
rect 16078 9220 16084 9222
rect 15776 9200 16084 9220
rect 15776 8188 16084 8208
rect 15776 8186 15782 8188
rect 15838 8186 15862 8188
rect 15918 8186 15942 8188
rect 15998 8186 16022 8188
rect 16078 8186 16084 8188
rect 15838 8134 15840 8186
rect 16020 8134 16022 8186
rect 15776 8132 15782 8134
rect 15838 8132 15862 8134
rect 15918 8132 15942 8134
rect 15998 8132 16022 8134
rect 16078 8132 16084 8134
rect 15776 8112 16084 8132
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 15776 7100 16084 7120
rect 15776 7098 15782 7100
rect 15838 7098 15862 7100
rect 15918 7098 15942 7100
rect 15998 7098 16022 7100
rect 16078 7098 16084 7100
rect 15838 7046 15840 7098
rect 16020 7046 16022 7098
rect 15776 7044 15782 7046
rect 15838 7044 15862 7046
rect 15918 7044 15942 7046
rect 15998 7044 16022 7046
rect 16078 7044 16084 7046
rect 15776 7024 16084 7044
rect 16224 6662 16252 7142
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15580 5914 15608 6258
rect 15776 6012 16084 6032
rect 15776 6010 15782 6012
rect 15838 6010 15862 6012
rect 15918 6010 15942 6012
rect 15998 6010 16022 6012
rect 16078 6010 16084 6012
rect 15838 5958 15840 6010
rect 16020 5958 16022 6010
rect 15776 5956 15782 5958
rect 15838 5956 15862 5958
rect 15918 5956 15942 5958
rect 15998 5956 16022 5958
rect 16078 5956 16084 5958
rect 15776 5936 16084 5956
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 16224 5710 16252 6598
rect 16776 5914 16804 6666
rect 17512 6322 17540 9658
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16960 5710 16988 6054
rect 17328 5914 17356 6258
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 15568 5568 15620 5574
rect 17880 5545 17908 5646
rect 15568 5510 15620 5516
rect 17866 5536 17922 5545
rect 15580 4622 15608 5510
rect 17866 5471 17922 5480
rect 15776 4924 16084 4944
rect 15776 4922 15782 4924
rect 15838 4922 15862 4924
rect 15918 4922 15942 4924
rect 15998 4922 16022 4924
rect 16078 4922 16084 4924
rect 15838 4870 15840 4922
rect 16020 4870 16022 4922
rect 15776 4868 15782 4870
rect 15838 4868 15862 4870
rect 15918 4868 15942 4870
rect 15998 4868 16022 4870
rect 16078 4868 16084 4870
rect 15776 4848 16084 4868
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 15776 3836 16084 3856
rect 15776 3834 15782 3836
rect 15838 3834 15862 3836
rect 15918 3834 15942 3836
rect 15998 3834 16022 3836
rect 16078 3834 16084 3836
rect 15838 3782 15840 3834
rect 16020 3782 16022 3834
rect 15776 3780 15782 3782
rect 15838 3780 15862 3782
rect 15918 3780 15942 3782
rect 15998 3780 16022 3782
rect 16078 3780 16084 3782
rect 15776 3760 16084 3780
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 6880 3292 7188 3312
rect 6880 3290 6886 3292
rect 6942 3290 6966 3292
rect 7022 3290 7046 3292
rect 7102 3290 7126 3292
rect 7182 3290 7188 3292
rect 6942 3238 6944 3290
rect 7124 3238 7126 3290
rect 6880 3236 6886 3238
rect 6942 3236 6966 3238
rect 7022 3236 7046 3238
rect 7102 3236 7126 3238
rect 7182 3236 7188 3238
rect 6880 3216 7188 3236
rect 3915 2748 4223 2768
rect 3915 2746 3921 2748
rect 3977 2746 4001 2748
rect 4057 2746 4081 2748
rect 4137 2746 4161 2748
rect 4217 2746 4223 2748
rect 3977 2694 3979 2746
rect 4159 2694 4161 2746
rect 3915 2692 3921 2694
rect 3977 2692 4001 2694
rect 4057 2692 4081 2694
rect 4137 2692 4161 2694
rect 4217 2692 4223 2694
rect 3915 2672 4223 2692
rect 9140 2650 9168 3470
rect 12811 3292 13119 3312
rect 12811 3290 12817 3292
rect 12873 3290 12897 3292
rect 12953 3290 12977 3292
rect 13033 3290 13057 3292
rect 13113 3290 13119 3292
rect 12873 3238 12875 3290
rect 13055 3238 13057 3290
rect 12811 3236 12817 3238
rect 12873 3236 12897 3238
rect 12953 3236 12977 3238
rect 13033 3236 13057 3238
rect 13113 3236 13119 3238
rect 12811 3216 13119 3236
rect 9846 2748 10154 2768
rect 9846 2746 9852 2748
rect 9908 2746 9932 2748
rect 9988 2746 10012 2748
rect 10068 2746 10092 2748
rect 10148 2746 10154 2748
rect 9908 2694 9910 2746
rect 10090 2694 10092 2746
rect 9846 2692 9852 2694
rect 9908 2692 9932 2694
rect 9988 2692 10012 2694
rect 10068 2692 10092 2694
rect 10148 2692 10154 2694
rect 9846 2672 10154 2692
rect 15776 2748 16084 2768
rect 15776 2746 15782 2748
rect 15838 2746 15862 2748
rect 15918 2746 15942 2748
rect 15998 2746 16022 2748
rect 16078 2746 16084 2748
rect 15838 2694 15840 2746
rect 16020 2694 16022 2746
rect 15776 2692 15782 2694
rect 15838 2692 15862 2694
rect 15918 2692 15942 2694
rect 15998 2692 16022 2694
rect 16078 2692 16084 2694
rect 15776 2672 16084 2692
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 16868 2446 16896 3878
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 32 800 60 2382
rect 6880 2204 7188 2224
rect 6880 2202 6886 2204
rect 6942 2202 6966 2204
rect 7022 2202 7046 2204
rect 7102 2202 7126 2204
rect 7182 2202 7188 2204
rect 6942 2150 6944 2202
rect 7124 2150 7126 2202
rect 6880 2148 6886 2150
rect 6942 2148 6966 2150
rect 7022 2148 7046 2150
rect 7102 2148 7126 2150
rect 7182 2148 7188 2150
rect 6880 2128 7188 2148
rect 8404 800 8432 2382
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 12811 2204 13119 2224
rect 12811 2202 12817 2204
rect 12873 2202 12897 2204
rect 12953 2202 12977 2204
rect 13033 2202 13057 2204
rect 13113 2202 13119 2204
rect 12873 2150 12875 2202
rect 13055 2150 13057 2202
rect 12811 2148 12817 2150
rect 12873 2148 12897 2150
rect 12953 2148 12977 2150
rect 13033 2148 13057 2150
rect 13113 2148 13119 2150
rect 12811 2128 13119 2148
rect 16776 800 16804 2246
rect 18 0 74 800
rect 8390 0 8446 800
rect 16762 0 16818 800
<< via2 >>
rect 3921 47354 3977 47356
rect 4001 47354 4057 47356
rect 4081 47354 4137 47356
rect 4161 47354 4217 47356
rect 3921 47302 3967 47354
rect 3967 47302 3977 47354
rect 4001 47302 4031 47354
rect 4031 47302 4043 47354
rect 4043 47302 4057 47354
rect 4081 47302 4095 47354
rect 4095 47302 4107 47354
rect 4107 47302 4137 47354
rect 4161 47302 4171 47354
rect 4171 47302 4217 47354
rect 3921 47300 3977 47302
rect 4001 47300 4057 47302
rect 4081 47300 4137 47302
rect 4161 47300 4217 47302
rect 9852 47354 9908 47356
rect 9932 47354 9988 47356
rect 10012 47354 10068 47356
rect 10092 47354 10148 47356
rect 9852 47302 9898 47354
rect 9898 47302 9908 47354
rect 9932 47302 9962 47354
rect 9962 47302 9974 47354
rect 9974 47302 9988 47354
rect 10012 47302 10026 47354
rect 10026 47302 10038 47354
rect 10038 47302 10068 47354
rect 10092 47302 10102 47354
rect 10102 47302 10148 47354
rect 9852 47300 9908 47302
rect 9932 47300 9988 47302
rect 10012 47300 10068 47302
rect 10092 47300 10148 47302
rect 15782 47354 15838 47356
rect 15862 47354 15918 47356
rect 15942 47354 15998 47356
rect 16022 47354 16078 47356
rect 15782 47302 15828 47354
rect 15828 47302 15838 47354
rect 15862 47302 15892 47354
rect 15892 47302 15904 47354
rect 15904 47302 15918 47354
rect 15942 47302 15956 47354
rect 15956 47302 15968 47354
rect 15968 47302 15998 47354
rect 16022 47302 16032 47354
rect 16032 47302 16078 47354
rect 15782 47300 15838 47302
rect 15862 47300 15918 47302
rect 15942 47300 15998 47302
rect 16022 47300 16078 47302
rect 1858 44240 1914 44296
rect 1398 35400 1454 35456
rect 1490 26560 1546 26616
rect 6886 46810 6942 46812
rect 6966 46810 7022 46812
rect 7046 46810 7102 46812
rect 7126 46810 7182 46812
rect 6886 46758 6932 46810
rect 6932 46758 6942 46810
rect 6966 46758 6996 46810
rect 6996 46758 7008 46810
rect 7008 46758 7022 46810
rect 7046 46758 7060 46810
rect 7060 46758 7072 46810
rect 7072 46758 7102 46810
rect 7126 46758 7136 46810
rect 7136 46758 7182 46810
rect 6886 46756 6942 46758
rect 6966 46756 7022 46758
rect 7046 46756 7102 46758
rect 7126 46756 7182 46758
rect 12817 46810 12873 46812
rect 12897 46810 12953 46812
rect 12977 46810 13033 46812
rect 13057 46810 13113 46812
rect 12817 46758 12863 46810
rect 12863 46758 12873 46810
rect 12897 46758 12927 46810
rect 12927 46758 12939 46810
rect 12939 46758 12953 46810
rect 12977 46758 12991 46810
rect 12991 46758 13003 46810
rect 13003 46758 13033 46810
rect 13057 46758 13067 46810
rect 13067 46758 13113 46810
rect 12817 46756 12873 46758
rect 12897 46756 12953 46758
rect 12977 46756 13033 46758
rect 13057 46756 13113 46758
rect 3921 46266 3977 46268
rect 4001 46266 4057 46268
rect 4081 46266 4137 46268
rect 4161 46266 4217 46268
rect 3921 46214 3967 46266
rect 3967 46214 3977 46266
rect 4001 46214 4031 46266
rect 4031 46214 4043 46266
rect 4043 46214 4057 46266
rect 4081 46214 4095 46266
rect 4095 46214 4107 46266
rect 4107 46214 4137 46266
rect 4161 46214 4171 46266
rect 4171 46214 4217 46266
rect 3921 46212 3977 46214
rect 4001 46212 4057 46214
rect 4081 46212 4137 46214
rect 4161 46212 4217 46214
rect 9852 46266 9908 46268
rect 9932 46266 9988 46268
rect 10012 46266 10068 46268
rect 10092 46266 10148 46268
rect 9852 46214 9898 46266
rect 9898 46214 9908 46266
rect 9932 46214 9962 46266
rect 9962 46214 9974 46266
rect 9974 46214 9988 46266
rect 10012 46214 10026 46266
rect 10026 46214 10038 46266
rect 10038 46214 10068 46266
rect 10092 46214 10102 46266
rect 10102 46214 10148 46266
rect 9852 46212 9908 46214
rect 9932 46212 9988 46214
rect 10012 46212 10068 46214
rect 10092 46212 10148 46214
rect 15782 46266 15838 46268
rect 15862 46266 15918 46268
rect 15942 46266 15998 46268
rect 16022 46266 16078 46268
rect 15782 46214 15828 46266
rect 15828 46214 15838 46266
rect 15862 46214 15892 46266
rect 15892 46214 15904 46266
rect 15904 46214 15918 46266
rect 15942 46214 15956 46266
rect 15956 46214 15968 46266
rect 15968 46214 15998 46266
rect 16022 46214 16032 46266
rect 16032 46214 16078 46266
rect 15782 46212 15838 46214
rect 15862 46212 15918 46214
rect 15942 46212 15998 46214
rect 16022 46212 16078 46214
rect 6886 45722 6942 45724
rect 6966 45722 7022 45724
rect 7046 45722 7102 45724
rect 7126 45722 7182 45724
rect 6886 45670 6932 45722
rect 6932 45670 6942 45722
rect 6966 45670 6996 45722
rect 6996 45670 7008 45722
rect 7008 45670 7022 45722
rect 7046 45670 7060 45722
rect 7060 45670 7072 45722
rect 7072 45670 7102 45722
rect 7126 45670 7136 45722
rect 7136 45670 7182 45722
rect 6886 45668 6942 45670
rect 6966 45668 7022 45670
rect 7046 45668 7102 45670
rect 7126 45668 7182 45670
rect 3921 45178 3977 45180
rect 4001 45178 4057 45180
rect 4081 45178 4137 45180
rect 4161 45178 4217 45180
rect 3921 45126 3967 45178
rect 3967 45126 3977 45178
rect 4001 45126 4031 45178
rect 4031 45126 4043 45178
rect 4043 45126 4057 45178
rect 4081 45126 4095 45178
rect 4095 45126 4107 45178
rect 4107 45126 4137 45178
rect 4161 45126 4171 45178
rect 4171 45126 4217 45178
rect 3921 45124 3977 45126
rect 4001 45124 4057 45126
rect 4081 45124 4137 45126
rect 4161 45124 4217 45126
rect 3921 44090 3977 44092
rect 4001 44090 4057 44092
rect 4081 44090 4137 44092
rect 4161 44090 4217 44092
rect 3921 44038 3967 44090
rect 3967 44038 3977 44090
rect 4001 44038 4031 44090
rect 4031 44038 4043 44090
rect 4043 44038 4057 44090
rect 4081 44038 4095 44090
rect 4095 44038 4107 44090
rect 4107 44038 4137 44090
rect 4161 44038 4171 44090
rect 4171 44038 4217 44090
rect 3921 44036 3977 44038
rect 4001 44036 4057 44038
rect 4081 44036 4137 44038
rect 4161 44036 4217 44038
rect 3921 43002 3977 43004
rect 4001 43002 4057 43004
rect 4081 43002 4137 43004
rect 4161 43002 4217 43004
rect 3921 42950 3967 43002
rect 3967 42950 3977 43002
rect 4001 42950 4031 43002
rect 4031 42950 4043 43002
rect 4043 42950 4057 43002
rect 4081 42950 4095 43002
rect 4095 42950 4107 43002
rect 4107 42950 4137 43002
rect 4161 42950 4171 43002
rect 4171 42950 4217 43002
rect 3921 42948 3977 42950
rect 4001 42948 4057 42950
rect 4081 42948 4137 42950
rect 4161 42948 4217 42950
rect 3921 41914 3977 41916
rect 4001 41914 4057 41916
rect 4081 41914 4137 41916
rect 4161 41914 4217 41916
rect 3921 41862 3967 41914
rect 3967 41862 3977 41914
rect 4001 41862 4031 41914
rect 4031 41862 4043 41914
rect 4043 41862 4057 41914
rect 4081 41862 4095 41914
rect 4095 41862 4107 41914
rect 4107 41862 4137 41914
rect 4161 41862 4171 41914
rect 4171 41862 4217 41914
rect 3921 41860 3977 41862
rect 4001 41860 4057 41862
rect 4081 41860 4137 41862
rect 4161 41860 4217 41862
rect 3921 40826 3977 40828
rect 4001 40826 4057 40828
rect 4081 40826 4137 40828
rect 4161 40826 4217 40828
rect 3921 40774 3967 40826
rect 3967 40774 3977 40826
rect 4001 40774 4031 40826
rect 4031 40774 4043 40826
rect 4043 40774 4057 40826
rect 4081 40774 4095 40826
rect 4095 40774 4107 40826
rect 4107 40774 4137 40826
rect 4161 40774 4171 40826
rect 4171 40774 4217 40826
rect 3921 40772 3977 40774
rect 4001 40772 4057 40774
rect 4081 40772 4137 40774
rect 4161 40772 4217 40774
rect 3921 39738 3977 39740
rect 4001 39738 4057 39740
rect 4081 39738 4137 39740
rect 4161 39738 4217 39740
rect 3921 39686 3967 39738
rect 3967 39686 3977 39738
rect 4001 39686 4031 39738
rect 4031 39686 4043 39738
rect 4043 39686 4057 39738
rect 4081 39686 4095 39738
rect 4095 39686 4107 39738
rect 4107 39686 4137 39738
rect 4161 39686 4171 39738
rect 4171 39686 4217 39738
rect 3921 39684 3977 39686
rect 4001 39684 4057 39686
rect 4081 39684 4137 39686
rect 4161 39684 4217 39686
rect 3921 38650 3977 38652
rect 4001 38650 4057 38652
rect 4081 38650 4137 38652
rect 4161 38650 4217 38652
rect 3921 38598 3967 38650
rect 3967 38598 3977 38650
rect 4001 38598 4031 38650
rect 4031 38598 4043 38650
rect 4043 38598 4057 38650
rect 4081 38598 4095 38650
rect 4095 38598 4107 38650
rect 4107 38598 4137 38650
rect 4161 38598 4171 38650
rect 4171 38598 4217 38650
rect 3921 38596 3977 38598
rect 4001 38596 4057 38598
rect 4081 38596 4137 38598
rect 4161 38596 4217 38598
rect 3921 37562 3977 37564
rect 4001 37562 4057 37564
rect 4081 37562 4137 37564
rect 4161 37562 4217 37564
rect 3921 37510 3967 37562
rect 3967 37510 3977 37562
rect 4001 37510 4031 37562
rect 4031 37510 4043 37562
rect 4043 37510 4057 37562
rect 4081 37510 4095 37562
rect 4095 37510 4107 37562
rect 4107 37510 4137 37562
rect 4161 37510 4171 37562
rect 4171 37510 4217 37562
rect 3921 37508 3977 37510
rect 4001 37508 4057 37510
rect 4081 37508 4137 37510
rect 4161 37508 4217 37510
rect 3921 36474 3977 36476
rect 4001 36474 4057 36476
rect 4081 36474 4137 36476
rect 4161 36474 4217 36476
rect 3921 36422 3967 36474
rect 3967 36422 3977 36474
rect 4001 36422 4031 36474
rect 4031 36422 4043 36474
rect 4043 36422 4057 36474
rect 4081 36422 4095 36474
rect 4095 36422 4107 36474
rect 4107 36422 4137 36474
rect 4161 36422 4171 36474
rect 4171 36422 4217 36474
rect 3921 36420 3977 36422
rect 4001 36420 4057 36422
rect 4081 36420 4137 36422
rect 4161 36420 4217 36422
rect 3921 35386 3977 35388
rect 4001 35386 4057 35388
rect 4081 35386 4137 35388
rect 4161 35386 4217 35388
rect 3921 35334 3967 35386
rect 3967 35334 3977 35386
rect 4001 35334 4031 35386
rect 4031 35334 4043 35386
rect 4043 35334 4057 35386
rect 4081 35334 4095 35386
rect 4095 35334 4107 35386
rect 4107 35334 4137 35386
rect 4161 35334 4171 35386
rect 4171 35334 4217 35386
rect 3921 35332 3977 35334
rect 4001 35332 4057 35334
rect 4081 35332 4137 35334
rect 4161 35332 4217 35334
rect 6886 44634 6942 44636
rect 6966 44634 7022 44636
rect 7046 44634 7102 44636
rect 7126 44634 7182 44636
rect 6886 44582 6932 44634
rect 6932 44582 6942 44634
rect 6966 44582 6996 44634
rect 6996 44582 7008 44634
rect 7008 44582 7022 44634
rect 7046 44582 7060 44634
rect 7060 44582 7072 44634
rect 7072 44582 7102 44634
rect 7126 44582 7136 44634
rect 7136 44582 7182 44634
rect 6886 44580 6942 44582
rect 6966 44580 7022 44582
rect 7046 44580 7102 44582
rect 7126 44580 7182 44582
rect 6886 43546 6942 43548
rect 6966 43546 7022 43548
rect 7046 43546 7102 43548
rect 7126 43546 7182 43548
rect 6886 43494 6932 43546
rect 6932 43494 6942 43546
rect 6966 43494 6996 43546
rect 6996 43494 7008 43546
rect 7008 43494 7022 43546
rect 7046 43494 7060 43546
rect 7060 43494 7072 43546
rect 7072 43494 7102 43546
rect 7126 43494 7136 43546
rect 7136 43494 7182 43546
rect 6886 43492 6942 43494
rect 6966 43492 7022 43494
rect 7046 43492 7102 43494
rect 7126 43492 7182 43494
rect 6886 42458 6942 42460
rect 6966 42458 7022 42460
rect 7046 42458 7102 42460
rect 7126 42458 7182 42460
rect 6886 42406 6932 42458
rect 6932 42406 6942 42458
rect 6966 42406 6996 42458
rect 6996 42406 7008 42458
rect 7008 42406 7022 42458
rect 7046 42406 7060 42458
rect 7060 42406 7072 42458
rect 7072 42406 7102 42458
rect 7126 42406 7136 42458
rect 7136 42406 7182 42458
rect 6886 42404 6942 42406
rect 6966 42404 7022 42406
rect 7046 42404 7102 42406
rect 7126 42404 7182 42406
rect 6886 41370 6942 41372
rect 6966 41370 7022 41372
rect 7046 41370 7102 41372
rect 7126 41370 7182 41372
rect 6886 41318 6932 41370
rect 6932 41318 6942 41370
rect 6966 41318 6996 41370
rect 6996 41318 7008 41370
rect 7008 41318 7022 41370
rect 7046 41318 7060 41370
rect 7060 41318 7072 41370
rect 7072 41318 7102 41370
rect 7126 41318 7136 41370
rect 7136 41318 7182 41370
rect 6886 41316 6942 41318
rect 6966 41316 7022 41318
rect 7046 41316 7102 41318
rect 7126 41316 7182 41318
rect 6886 40282 6942 40284
rect 6966 40282 7022 40284
rect 7046 40282 7102 40284
rect 7126 40282 7182 40284
rect 6886 40230 6932 40282
rect 6932 40230 6942 40282
rect 6966 40230 6996 40282
rect 6996 40230 7008 40282
rect 7008 40230 7022 40282
rect 7046 40230 7060 40282
rect 7060 40230 7072 40282
rect 7072 40230 7102 40282
rect 7126 40230 7136 40282
rect 7136 40230 7182 40282
rect 6886 40228 6942 40230
rect 6966 40228 7022 40230
rect 7046 40228 7102 40230
rect 7126 40228 7182 40230
rect 6886 39194 6942 39196
rect 6966 39194 7022 39196
rect 7046 39194 7102 39196
rect 7126 39194 7182 39196
rect 6886 39142 6932 39194
rect 6932 39142 6942 39194
rect 6966 39142 6996 39194
rect 6996 39142 7008 39194
rect 7008 39142 7022 39194
rect 7046 39142 7060 39194
rect 7060 39142 7072 39194
rect 7072 39142 7102 39194
rect 7126 39142 7136 39194
rect 7136 39142 7182 39194
rect 6886 39140 6942 39142
rect 6966 39140 7022 39142
rect 7046 39140 7102 39142
rect 7126 39140 7182 39142
rect 3921 34298 3977 34300
rect 4001 34298 4057 34300
rect 4081 34298 4137 34300
rect 4161 34298 4217 34300
rect 3921 34246 3967 34298
rect 3967 34246 3977 34298
rect 4001 34246 4031 34298
rect 4031 34246 4043 34298
rect 4043 34246 4057 34298
rect 4081 34246 4095 34298
rect 4095 34246 4107 34298
rect 4107 34246 4137 34298
rect 4161 34246 4171 34298
rect 4171 34246 4217 34298
rect 3921 34244 3977 34246
rect 4001 34244 4057 34246
rect 4081 34244 4137 34246
rect 4161 34244 4217 34246
rect 3921 33210 3977 33212
rect 4001 33210 4057 33212
rect 4081 33210 4137 33212
rect 4161 33210 4217 33212
rect 3921 33158 3967 33210
rect 3967 33158 3977 33210
rect 4001 33158 4031 33210
rect 4031 33158 4043 33210
rect 4043 33158 4057 33210
rect 4081 33158 4095 33210
rect 4095 33158 4107 33210
rect 4107 33158 4137 33210
rect 4161 33158 4171 33210
rect 4171 33158 4217 33210
rect 3921 33156 3977 33158
rect 4001 33156 4057 33158
rect 4081 33156 4137 33158
rect 4161 33156 4217 33158
rect 3921 32122 3977 32124
rect 4001 32122 4057 32124
rect 4081 32122 4137 32124
rect 4161 32122 4217 32124
rect 3921 32070 3967 32122
rect 3967 32070 3977 32122
rect 4001 32070 4031 32122
rect 4031 32070 4043 32122
rect 4043 32070 4057 32122
rect 4081 32070 4095 32122
rect 4095 32070 4107 32122
rect 4107 32070 4137 32122
rect 4161 32070 4171 32122
rect 4171 32070 4217 32122
rect 3921 32068 3977 32070
rect 4001 32068 4057 32070
rect 4081 32068 4137 32070
rect 4161 32068 4217 32070
rect 3921 31034 3977 31036
rect 4001 31034 4057 31036
rect 4081 31034 4137 31036
rect 4161 31034 4217 31036
rect 3921 30982 3967 31034
rect 3967 30982 3977 31034
rect 4001 30982 4031 31034
rect 4031 30982 4043 31034
rect 4043 30982 4057 31034
rect 4081 30982 4095 31034
rect 4095 30982 4107 31034
rect 4107 30982 4137 31034
rect 4161 30982 4171 31034
rect 4171 30982 4217 31034
rect 3921 30980 3977 30982
rect 4001 30980 4057 30982
rect 4081 30980 4137 30982
rect 4161 30980 4217 30982
rect 3921 29946 3977 29948
rect 4001 29946 4057 29948
rect 4081 29946 4137 29948
rect 4161 29946 4217 29948
rect 3921 29894 3967 29946
rect 3967 29894 3977 29946
rect 4001 29894 4031 29946
rect 4031 29894 4043 29946
rect 4043 29894 4057 29946
rect 4081 29894 4095 29946
rect 4095 29894 4107 29946
rect 4107 29894 4137 29946
rect 4161 29894 4171 29946
rect 4171 29894 4217 29946
rect 3921 29892 3977 29894
rect 4001 29892 4057 29894
rect 4081 29892 4137 29894
rect 4161 29892 4217 29894
rect 3921 28858 3977 28860
rect 4001 28858 4057 28860
rect 4081 28858 4137 28860
rect 4161 28858 4217 28860
rect 3921 28806 3967 28858
rect 3967 28806 3977 28858
rect 4001 28806 4031 28858
rect 4031 28806 4043 28858
rect 4043 28806 4057 28858
rect 4081 28806 4095 28858
rect 4095 28806 4107 28858
rect 4107 28806 4137 28858
rect 4161 28806 4171 28858
rect 4171 28806 4217 28858
rect 3921 28804 3977 28806
rect 4001 28804 4057 28806
rect 4081 28804 4137 28806
rect 4161 28804 4217 28806
rect 3921 27770 3977 27772
rect 4001 27770 4057 27772
rect 4081 27770 4137 27772
rect 4161 27770 4217 27772
rect 3921 27718 3967 27770
rect 3967 27718 3977 27770
rect 4001 27718 4031 27770
rect 4031 27718 4043 27770
rect 4043 27718 4057 27770
rect 4081 27718 4095 27770
rect 4095 27718 4107 27770
rect 4107 27718 4137 27770
rect 4161 27718 4171 27770
rect 4171 27718 4217 27770
rect 3921 27716 3977 27718
rect 4001 27716 4057 27718
rect 4081 27716 4137 27718
rect 4161 27716 4217 27718
rect 3921 26682 3977 26684
rect 4001 26682 4057 26684
rect 4081 26682 4137 26684
rect 4161 26682 4217 26684
rect 3921 26630 3967 26682
rect 3967 26630 3977 26682
rect 4001 26630 4031 26682
rect 4031 26630 4043 26682
rect 4043 26630 4057 26682
rect 4081 26630 4095 26682
rect 4095 26630 4107 26682
rect 4107 26630 4137 26682
rect 4161 26630 4171 26682
rect 4171 26630 4217 26682
rect 3921 26628 3977 26630
rect 4001 26628 4057 26630
rect 4081 26628 4137 26630
rect 4161 26628 4217 26630
rect 3921 25594 3977 25596
rect 4001 25594 4057 25596
rect 4081 25594 4137 25596
rect 4161 25594 4217 25596
rect 3921 25542 3967 25594
rect 3967 25542 3977 25594
rect 4001 25542 4031 25594
rect 4031 25542 4043 25594
rect 4043 25542 4057 25594
rect 4081 25542 4095 25594
rect 4095 25542 4107 25594
rect 4107 25542 4137 25594
rect 4161 25542 4171 25594
rect 4171 25542 4217 25594
rect 3921 25540 3977 25542
rect 4001 25540 4057 25542
rect 4081 25540 4137 25542
rect 4161 25540 4217 25542
rect 3921 24506 3977 24508
rect 4001 24506 4057 24508
rect 4081 24506 4137 24508
rect 4161 24506 4217 24508
rect 3921 24454 3967 24506
rect 3967 24454 3977 24506
rect 4001 24454 4031 24506
rect 4031 24454 4043 24506
rect 4043 24454 4057 24506
rect 4081 24454 4095 24506
rect 4095 24454 4107 24506
rect 4107 24454 4137 24506
rect 4161 24454 4171 24506
rect 4171 24454 4217 24506
rect 3921 24452 3977 24454
rect 4001 24452 4057 24454
rect 4081 24452 4137 24454
rect 4161 24452 4217 24454
rect 6886 38106 6942 38108
rect 6966 38106 7022 38108
rect 7046 38106 7102 38108
rect 7126 38106 7182 38108
rect 6886 38054 6932 38106
rect 6932 38054 6942 38106
rect 6966 38054 6996 38106
rect 6996 38054 7008 38106
rect 7008 38054 7022 38106
rect 7046 38054 7060 38106
rect 7060 38054 7072 38106
rect 7072 38054 7102 38106
rect 7126 38054 7136 38106
rect 7136 38054 7182 38106
rect 6886 38052 6942 38054
rect 6966 38052 7022 38054
rect 7046 38052 7102 38054
rect 7126 38052 7182 38054
rect 6886 37018 6942 37020
rect 6966 37018 7022 37020
rect 7046 37018 7102 37020
rect 7126 37018 7182 37020
rect 6886 36966 6932 37018
rect 6932 36966 6942 37018
rect 6966 36966 6996 37018
rect 6996 36966 7008 37018
rect 7008 36966 7022 37018
rect 7046 36966 7060 37018
rect 7060 36966 7072 37018
rect 7072 36966 7102 37018
rect 7126 36966 7136 37018
rect 7136 36966 7182 37018
rect 6886 36964 6942 36966
rect 6966 36964 7022 36966
rect 7046 36964 7102 36966
rect 7126 36964 7182 36966
rect 6886 35930 6942 35932
rect 6966 35930 7022 35932
rect 7046 35930 7102 35932
rect 7126 35930 7182 35932
rect 6886 35878 6932 35930
rect 6932 35878 6942 35930
rect 6966 35878 6996 35930
rect 6996 35878 7008 35930
rect 7008 35878 7022 35930
rect 7046 35878 7060 35930
rect 7060 35878 7072 35930
rect 7072 35878 7102 35930
rect 7126 35878 7136 35930
rect 7136 35878 7182 35930
rect 6886 35876 6942 35878
rect 6966 35876 7022 35878
rect 7046 35876 7102 35878
rect 7126 35876 7182 35878
rect 6886 34842 6942 34844
rect 6966 34842 7022 34844
rect 7046 34842 7102 34844
rect 7126 34842 7182 34844
rect 6886 34790 6932 34842
rect 6932 34790 6942 34842
rect 6966 34790 6996 34842
rect 6996 34790 7008 34842
rect 7008 34790 7022 34842
rect 7046 34790 7060 34842
rect 7060 34790 7072 34842
rect 7072 34790 7102 34842
rect 7126 34790 7136 34842
rect 7136 34790 7182 34842
rect 6886 34788 6942 34790
rect 6966 34788 7022 34790
rect 7046 34788 7102 34790
rect 7126 34788 7182 34790
rect 5998 33088 6054 33144
rect 3921 23418 3977 23420
rect 4001 23418 4057 23420
rect 4081 23418 4137 23420
rect 4161 23418 4217 23420
rect 3921 23366 3967 23418
rect 3967 23366 3977 23418
rect 4001 23366 4031 23418
rect 4031 23366 4043 23418
rect 4043 23366 4057 23418
rect 4081 23366 4095 23418
rect 4095 23366 4107 23418
rect 4107 23366 4137 23418
rect 4161 23366 4171 23418
rect 4171 23366 4217 23418
rect 3921 23364 3977 23366
rect 4001 23364 4057 23366
rect 4081 23364 4137 23366
rect 4161 23364 4217 23366
rect 3921 22330 3977 22332
rect 4001 22330 4057 22332
rect 4081 22330 4137 22332
rect 4161 22330 4217 22332
rect 3921 22278 3967 22330
rect 3967 22278 3977 22330
rect 4001 22278 4031 22330
rect 4031 22278 4043 22330
rect 4043 22278 4057 22330
rect 4081 22278 4095 22330
rect 4095 22278 4107 22330
rect 4107 22278 4137 22330
rect 4161 22278 4171 22330
rect 4171 22278 4217 22330
rect 3921 22276 3977 22278
rect 4001 22276 4057 22278
rect 4081 22276 4137 22278
rect 4161 22276 4217 22278
rect 1398 17720 1454 17776
rect 3921 21242 3977 21244
rect 4001 21242 4057 21244
rect 4081 21242 4137 21244
rect 4161 21242 4217 21244
rect 3921 21190 3967 21242
rect 3967 21190 3977 21242
rect 4001 21190 4031 21242
rect 4031 21190 4043 21242
rect 4043 21190 4057 21242
rect 4081 21190 4095 21242
rect 4095 21190 4107 21242
rect 4107 21190 4137 21242
rect 4161 21190 4171 21242
rect 4171 21190 4217 21242
rect 3921 21188 3977 21190
rect 4001 21188 4057 21190
rect 4081 21188 4137 21190
rect 4161 21188 4217 21190
rect 3921 20154 3977 20156
rect 4001 20154 4057 20156
rect 4081 20154 4137 20156
rect 4161 20154 4217 20156
rect 3921 20102 3967 20154
rect 3967 20102 3977 20154
rect 4001 20102 4031 20154
rect 4031 20102 4043 20154
rect 4043 20102 4057 20154
rect 4081 20102 4095 20154
rect 4095 20102 4107 20154
rect 4107 20102 4137 20154
rect 4161 20102 4171 20154
rect 4171 20102 4217 20154
rect 3921 20100 3977 20102
rect 4001 20100 4057 20102
rect 4081 20100 4137 20102
rect 4161 20100 4217 20102
rect 3921 19066 3977 19068
rect 4001 19066 4057 19068
rect 4081 19066 4137 19068
rect 4161 19066 4217 19068
rect 3921 19014 3967 19066
rect 3967 19014 3977 19066
rect 4001 19014 4031 19066
rect 4031 19014 4043 19066
rect 4043 19014 4057 19066
rect 4081 19014 4095 19066
rect 4095 19014 4107 19066
rect 4107 19014 4137 19066
rect 4161 19014 4171 19066
rect 4171 19014 4217 19066
rect 3921 19012 3977 19014
rect 4001 19012 4057 19014
rect 4081 19012 4137 19014
rect 4161 19012 4217 19014
rect 3921 17978 3977 17980
rect 4001 17978 4057 17980
rect 4081 17978 4137 17980
rect 4161 17978 4217 17980
rect 3921 17926 3967 17978
rect 3967 17926 3977 17978
rect 4001 17926 4031 17978
rect 4031 17926 4043 17978
rect 4043 17926 4057 17978
rect 4081 17926 4095 17978
rect 4095 17926 4107 17978
rect 4107 17926 4137 17978
rect 4161 17926 4171 17978
rect 4171 17926 4217 17978
rect 3921 17924 3977 17926
rect 4001 17924 4057 17926
rect 4081 17924 4137 17926
rect 4161 17924 4217 17926
rect 3921 16890 3977 16892
rect 4001 16890 4057 16892
rect 4081 16890 4137 16892
rect 4161 16890 4217 16892
rect 3921 16838 3967 16890
rect 3967 16838 3977 16890
rect 4001 16838 4031 16890
rect 4031 16838 4043 16890
rect 4043 16838 4057 16890
rect 4081 16838 4095 16890
rect 4095 16838 4107 16890
rect 4107 16838 4137 16890
rect 4161 16838 4171 16890
rect 4171 16838 4217 16890
rect 3921 16836 3977 16838
rect 4001 16836 4057 16838
rect 4081 16836 4137 16838
rect 4161 16836 4217 16838
rect 3921 15802 3977 15804
rect 4001 15802 4057 15804
rect 4081 15802 4137 15804
rect 4161 15802 4217 15804
rect 3921 15750 3967 15802
rect 3967 15750 3977 15802
rect 4001 15750 4031 15802
rect 4031 15750 4043 15802
rect 4043 15750 4057 15802
rect 4081 15750 4095 15802
rect 4095 15750 4107 15802
rect 4107 15750 4137 15802
rect 4161 15750 4171 15802
rect 4171 15750 4217 15802
rect 3921 15748 3977 15750
rect 4001 15748 4057 15750
rect 4081 15748 4137 15750
rect 4161 15748 4217 15750
rect 3921 14714 3977 14716
rect 4001 14714 4057 14716
rect 4081 14714 4137 14716
rect 4161 14714 4217 14716
rect 3921 14662 3967 14714
rect 3967 14662 3977 14714
rect 4001 14662 4031 14714
rect 4031 14662 4043 14714
rect 4043 14662 4057 14714
rect 4081 14662 4095 14714
rect 4095 14662 4107 14714
rect 4107 14662 4137 14714
rect 4161 14662 4171 14714
rect 4171 14662 4217 14714
rect 3921 14660 3977 14662
rect 4001 14660 4057 14662
rect 4081 14660 4137 14662
rect 4161 14660 4217 14662
rect 6886 33754 6942 33756
rect 6966 33754 7022 33756
rect 7046 33754 7102 33756
rect 7126 33754 7182 33756
rect 6886 33702 6932 33754
rect 6932 33702 6942 33754
rect 6966 33702 6996 33754
rect 6996 33702 7008 33754
rect 7008 33702 7022 33754
rect 7046 33702 7060 33754
rect 7060 33702 7072 33754
rect 7072 33702 7102 33754
rect 7126 33702 7136 33754
rect 7136 33702 7182 33754
rect 6886 33700 6942 33702
rect 6966 33700 7022 33702
rect 7046 33700 7102 33702
rect 7126 33700 7182 33702
rect 6886 32666 6942 32668
rect 6966 32666 7022 32668
rect 7046 32666 7102 32668
rect 7126 32666 7182 32668
rect 6886 32614 6932 32666
rect 6932 32614 6942 32666
rect 6966 32614 6996 32666
rect 6996 32614 7008 32666
rect 7008 32614 7022 32666
rect 7046 32614 7060 32666
rect 7060 32614 7072 32666
rect 7072 32614 7102 32666
rect 7126 32614 7136 32666
rect 7136 32614 7182 32666
rect 6886 32612 6942 32614
rect 6966 32612 7022 32614
rect 7046 32612 7102 32614
rect 7126 32612 7182 32614
rect 6886 31578 6942 31580
rect 6966 31578 7022 31580
rect 7046 31578 7102 31580
rect 7126 31578 7182 31580
rect 6886 31526 6932 31578
rect 6932 31526 6942 31578
rect 6966 31526 6996 31578
rect 6996 31526 7008 31578
rect 7008 31526 7022 31578
rect 7046 31526 7060 31578
rect 7060 31526 7072 31578
rect 7072 31526 7102 31578
rect 7126 31526 7136 31578
rect 7136 31526 7182 31578
rect 6886 31524 6942 31526
rect 6966 31524 7022 31526
rect 7046 31524 7102 31526
rect 7126 31524 7182 31526
rect 6886 30490 6942 30492
rect 6966 30490 7022 30492
rect 7046 30490 7102 30492
rect 7126 30490 7182 30492
rect 6886 30438 6932 30490
rect 6932 30438 6942 30490
rect 6966 30438 6996 30490
rect 6996 30438 7008 30490
rect 7008 30438 7022 30490
rect 7046 30438 7060 30490
rect 7060 30438 7072 30490
rect 7072 30438 7102 30490
rect 7126 30438 7136 30490
rect 7136 30438 7182 30490
rect 6886 30436 6942 30438
rect 6966 30436 7022 30438
rect 7046 30436 7102 30438
rect 7126 30436 7182 30438
rect 6886 29402 6942 29404
rect 6966 29402 7022 29404
rect 7046 29402 7102 29404
rect 7126 29402 7182 29404
rect 6886 29350 6932 29402
rect 6932 29350 6942 29402
rect 6966 29350 6996 29402
rect 6996 29350 7008 29402
rect 7008 29350 7022 29402
rect 7046 29350 7060 29402
rect 7060 29350 7072 29402
rect 7072 29350 7102 29402
rect 7126 29350 7136 29402
rect 7136 29350 7182 29402
rect 6886 29348 6942 29350
rect 6966 29348 7022 29350
rect 7046 29348 7102 29350
rect 7126 29348 7182 29350
rect 6886 28314 6942 28316
rect 6966 28314 7022 28316
rect 7046 28314 7102 28316
rect 7126 28314 7182 28316
rect 6886 28262 6932 28314
rect 6932 28262 6942 28314
rect 6966 28262 6996 28314
rect 6996 28262 7008 28314
rect 7008 28262 7022 28314
rect 7046 28262 7060 28314
rect 7060 28262 7072 28314
rect 7072 28262 7102 28314
rect 7126 28262 7136 28314
rect 7136 28262 7182 28314
rect 6886 28260 6942 28262
rect 6966 28260 7022 28262
rect 7046 28260 7102 28262
rect 7126 28260 7182 28262
rect 6886 27226 6942 27228
rect 6966 27226 7022 27228
rect 7046 27226 7102 27228
rect 7126 27226 7182 27228
rect 6886 27174 6932 27226
rect 6932 27174 6942 27226
rect 6966 27174 6996 27226
rect 6996 27174 7008 27226
rect 7008 27174 7022 27226
rect 7046 27174 7060 27226
rect 7060 27174 7072 27226
rect 7072 27174 7102 27226
rect 7126 27174 7136 27226
rect 7136 27174 7182 27226
rect 6886 27172 6942 27174
rect 6966 27172 7022 27174
rect 7046 27172 7102 27174
rect 7126 27172 7182 27174
rect 6886 26138 6942 26140
rect 6966 26138 7022 26140
rect 7046 26138 7102 26140
rect 7126 26138 7182 26140
rect 6886 26086 6932 26138
rect 6932 26086 6942 26138
rect 6966 26086 6996 26138
rect 6996 26086 7008 26138
rect 7008 26086 7022 26138
rect 7046 26086 7060 26138
rect 7060 26086 7072 26138
rect 7072 26086 7102 26138
rect 7126 26086 7136 26138
rect 7136 26086 7182 26138
rect 6886 26084 6942 26086
rect 6966 26084 7022 26086
rect 7046 26084 7102 26086
rect 7126 26084 7182 26086
rect 6886 25050 6942 25052
rect 6966 25050 7022 25052
rect 7046 25050 7102 25052
rect 7126 25050 7182 25052
rect 6886 24998 6932 25050
rect 6932 24998 6942 25050
rect 6966 24998 6996 25050
rect 6996 24998 7008 25050
rect 7008 24998 7022 25050
rect 7046 24998 7060 25050
rect 7060 24998 7072 25050
rect 7072 24998 7102 25050
rect 7126 24998 7136 25050
rect 7136 24998 7182 25050
rect 6886 24996 6942 24998
rect 6966 24996 7022 24998
rect 7046 24996 7102 24998
rect 7126 24996 7182 24998
rect 6886 23962 6942 23964
rect 6966 23962 7022 23964
rect 7046 23962 7102 23964
rect 7126 23962 7182 23964
rect 6886 23910 6932 23962
rect 6932 23910 6942 23962
rect 6966 23910 6996 23962
rect 6996 23910 7008 23962
rect 7008 23910 7022 23962
rect 7046 23910 7060 23962
rect 7060 23910 7072 23962
rect 7072 23910 7102 23962
rect 7126 23910 7136 23962
rect 7136 23910 7182 23962
rect 6886 23908 6942 23910
rect 6966 23908 7022 23910
rect 7046 23908 7102 23910
rect 7126 23908 7182 23910
rect 6886 22874 6942 22876
rect 6966 22874 7022 22876
rect 7046 22874 7102 22876
rect 7126 22874 7182 22876
rect 6886 22822 6932 22874
rect 6932 22822 6942 22874
rect 6966 22822 6996 22874
rect 6996 22822 7008 22874
rect 7008 22822 7022 22874
rect 7046 22822 7060 22874
rect 7060 22822 7072 22874
rect 7072 22822 7102 22874
rect 7126 22822 7136 22874
rect 7136 22822 7182 22874
rect 6886 22820 6942 22822
rect 6966 22820 7022 22822
rect 7046 22820 7102 22822
rect 7126 22820 7182 22822
rect 6886 21786 6942 21788
rect 6966 21786 7022 21788
rect 7046 21786 7102 21788
rect 7126 21786 7182 21788
rect 6886 21734 6932 21786
rect 6932 21734 6942 21786
rect 6966 21734 6996 21786
rect 6996 21734 7008 21786
rect 7008 21734 7022 21786
rect 7046 21734 7060 21786
rect 7060 21734 7072 21786
rect 7072 21734 7102 21786
rect 7126 21734 7136 21786
rect 7136 21734 7182 21786
rect 6886 21732 6942 21734
rect 6966 21732 7022 21734
rect 7046 21732 7102 21734
rect 7126 21732 7182 21734
rect 6886 20698 6942 20700
rect 6966 20698 7022 20700
rect 7046 20698 7102 20700
rect 7126 20698 7182 20700
rect 6886 20646 6932 20698
rect 6932 20646 6942 20698
rect 6966 20646 6996 20698
rect 6996 20646 7008 20698
rect 7008 20646 7022 20698
rect 7046 20646 7060 20698
rect 7060 20646 7072 20698
rect 7072 20646 7102 20698
rect 7126 20646 7136 20698
rect 7136 20646 7182 20698
rect 6886 20644 6942 20646
rect 6966 20644 7022 20646
rect 7046 20644 7102 20646
rect 7126 20644 7182 20646
rect 3921 13626 3977 13628
rect 4001 13626 4057 13628
rect 4081 13626 4137 13628
rect 4161 13626 4217 13628
rect 3921 13574 3967 13626
rect 3967 13574 3977 13626
rect 4001 13574 4031 13626
rect 4031 13574 4043 13626
rect 4043 13574 4057 13626
rect 4081 13574 4095 13626
rect 4095 13574 4107 13626
rect 4107 13574 4137 13626
rect 4161 13574 4171 13626
rect 4171 13574 4217 13626
rect 3921 13572 3977 13574
rect 4001 13572 4057 13574
rect 4081 13572 4137 13574
rect 4161 13572 4217 13574
rect 3921 12538 3977 12540
rect 4001 12538 4057 12540
rect 4081 12538 4137 12540
rect 4161 12538 4217 12540
rect 3921 12486 3967 12538
rect 3967 12486 3977 12538
rect 4001 12486 4031 12538
rect 4031 12486 4043 12538
rect 4043 12486 4057 12538
rect 4081 12486 4095 12538
rect 4095 12486 4107 12538
rect 4107 12486 4137 12538
rect 4161 12486 4171 12538
rect 4171 12486 4217 12538
rect 3921 12484 3977 12486
rect 4001 12484 4057 12486
rect 4081 12484 4137 12486
rect 4161 12484 4217 12486
rect 3921 11450 3977 11452
rect 4001 11450 4057 11452
rect 4081 11450 4137 11452
rect 4161 11450 4217 11452
rect 3921 11398 3967 11450
rect 3967 11398 3977 11450
rect 4001 11398 4031 11450
rect 4031 11398 4043 11450
rect 4043 11398 4057 11450
rect 4081 11398 4095 11450
rect 4095 11398 4107 11450
rect 4107 11398 4137 11450
rect 4161 11398 4171 11450
rect 4171 11398 4217 11450
rect 3921 11396 3977 11398
rect 4001 11396 4057 11398
rect 4081 11396 4137 11398
rect 4161 11396 4217 11398
rect 1398 8916 1400 8936
rect 1400 8916 1452 8936
rect 1452 8916 1454 8936
rect 1398 8880 1454 8916
rect 3921 10362 3977 10364
rect 4001 10362 4057 10364
rect 4081 10362 4137 10364
rect 4161 10362 4217 10364
rect 3921 10310 3967 10362
rect 3967 10310 3977 10362
rect 4001 10310 4031 10362
rect 4031 10310 4043 10362
rect 4043 10310 4057 10362
rect 4081 10310 4095 10362
rect 4095 10310 4107 10362
rect 4107 10310 4137 10362
rect 4161 10310 4171 10362
rect 4171 10310 4217 10362
rect 3921 10308 3977 10310
rect 4001 10308 4057 10310
rect 4081 10308 4137 10310
rect 4161 10308 4217 10310
rect 3921 9274 3977 9276
rect 4001 9274 4057 9276
rect 4081 9274 4137 9276
rect 4161 9274 4217 9276
rect 3921 9222 3967 9274
rect 3967 9222 3977 9274
rect 4001 9222 4031 9274
rect 4031 9222 4043 9274
rect 4043 9222 4057 9274
rect 4081 9222 4095 9274
rect 4095 9222 4107 9274
rect 4107 9222 4137 9274
rect 4161 9222 4171 9274
rect 4171 9222 4217 9274
rect 3921 9220 3977 9222
rect 4001 9220 4057 9222
rect 4081 9220 4137 9222
rect 4161 9220 4217 9222
rect 6886 19610 6942 19612
rect 6966 19610 7022 19612
rect 7046 19610 7102 19612
rect 7126 19610 7182 19612
rect 6886 19558 6932 19610
rect 6932 19558 6942 19610
rect 6966 19558 6996 19610
rect 6996 19558 7008 19610
rect 7008 19558 7022 19610
rect 7046 19558 7060 19610
rect 7060 19558 7072 19610
rect 7072 19558 7102 19610
rect 7126 19558 7136 19610
rect 7136 19558 7182 19610
rect 6886 19556 6942 19558
rect 6966 19556 7022 19558
rect 7046 19556 7102 19558
rect 7126 19556 7182 19558
rect 6886 18522 6942 18524
rect 6966 18522 7022 18524
rect 7046 18522 7102 18524
rect 7126 18522 7182 18524
rect 6886 18470 6932 18522
rect 6932 18470 6942 18522
rect 6966 18470 6996 18522
rect 6996 18470 7008 18522
rect 7008 18470 7022 18522
rect 7046 18470 7060 18522
rect 7060 18470 7072 18522
rect 7072 18470 7102 18522
rect 7126 18470 7136 18522
rect 7136 18470 7182 18522
rect 6886 18468 6942 18470
rect 6966 18468 7022 18470
rect 7046 18468 7102 18470
rect 7126 18468 7182 18470
rect 6090 15428 6146 15464
rect 6090 15408 6092 15428
rect 6092 15408 6144 15428
rect 6144 15408 6146 15428
rect 7930 33088 7986 33144
rect 12817 45722 12873 45724
rect 12897 45722 12953 45724
rect 12977 45722 13033 45724
rect 13057 45722 13113 45724
rect 12817 45670 12863 45722
rect 12863 45670 12873 45722
rect 12897 45670 12927 45722
rect 12927 45670 12939 45722
rect 12939 45670 12953 45722
rect 12977 45670 12991 45722
rect 12991 45670 13003 45722
rect 13003 45670 13033 45722
rect 13057 45670 13067 45722
rect 13067 45670 13113 45722
rect 12817 45668 12873 45670
rect 12897 45668 12953 45670
rect 12977 45668 13033 45670
rect 13057 45668 13113 45670
rect 9852 45178 9908 45180
rect 9932 45178 9988 45180
rect 10012 45178 10068 45180
rect 10092 45178 10148 45180
rect 9852 45126 9898 45178
rect 9898 45126 9908 45178
rect 9932 45126 9962 45178
rect 9962 45126 9974 45178
rect 9974 45126 9988 45178
rect 10012 45126 10026 45178
rect 10026 45126 10038 45178
rect 10038 45126 10068 45178
rect 10092 45126 10102 45178
rect 10102 45126 10148 45178
rect 9852 45124 9908 45126
rect 9932 45124 9988 45126
rect 10012 45124 10068 45126
rect 10092 45124 10148 45126
rect 9852 44090 9908 44092
rect 9932 44090 9988 44092
rect 10012 44090 10068 44092
rect 10092 44090 10148 44092
rect 9852 44038 9898 44090
rect 9898 44038 9908 44090
rect 9932 44038 9962 44090
rect 9962 44038 9974 44090
rect 9974 44038 9988 44090
rect 10012 44038 10026 44090
rect 10026 44038 10038 44090
rect 10038 44038 10068 44090
rect 10092 44038 10102 44090
rect 10102 44038 10148 44090
rect 9852 44036 9908 44038
rect 9932 44036 9988 44038
rect 10012 44036 10068 44038
rect 10092 44036 10148 44038
rect 9852 43002 9908 43004
rect 9932 43002 9988 43004
rect 10012 43002 10068 43004
rect 10092 43002 10148 43004
rect 9852 42950 9898 43002
rect 9898 42950 9908 43002
rect 9932 42950 9962 43002
rect 9962 42950 9974 43002
rect 9974 42950 9988 43002
rect 10012 42950 10026 43002
rect 10026 42950 10038 43002
rect 10038 42950 10068 43002
rect 10092 42950 10102 43002
rect 10102 42950 10148 43002
rect 9852 42948 9908 42950
rect 9932 42948 9988 42950
rect 10012 42948 10068 42950
rect 10092 42948 10148 42950
rect 9852 41914 9908 41916
rect 9932 41914 9988 41916
rect 10012 41914 10068 41916
rect 10092 41914 10148 41916
rect 9852 41862 9898 41914
rect 9898 41862 9908 41914
rect 9932 41862 9962 41914
rect 9962 41862 9974 41914
rect 9974 41862 9988 41914
rect 10012 41862 10026 41914
rect 10026 41862 10038 41914
rect 10038 41862 10068 41914
rect 10092 41862 10102 41914
rect 10102 41862 10148 41914
rect 9852 41860 9908 41862
rect 9932 41860 9988 41862
rect 10012 41860 10068 41862
rect 10092 41860 10148 41862
rect 9852 40826 9908 40828
rect 9932 40826 9988 40828
rect 10012 40826 10068 40828
rect 10092 40826 10148 40828
rect 9852 40774 9898 40826
rect 9898 40774 9908 40826
rect 9932 40774 9962 40826
rect 9962 40774 9974 40826
rect 9974 40774 9988 40826
rect 10012 40774 10026 40826
rect 10026 40774 10038 40826
rect 10038 40774 10068 40826
rect 10092 40774 10102 40826
rect 10102 40774 10148 40826
rect 9852 40772 9908 40774
rect 9932 40772 9988 40774
rect 10012 40772 10068 40774
rect 10092 40772 10148 40774
rect 9852 39738 9908 39740
rect 9932 39738 9988 39740
rect 10012 39738 10068 39740
rect 10092 39738 10148 39740
rect 9852 39686 9898 39738
rect 9898 39686 9908 39738
rect 9932 39686 9962 39738
rect 9962 39686 9974 39738
rect 9974 39686 9988 39738
rect 10012 39686 10026 39738
rect 10026 39686 10038 39738
rect 10038 39686 10068 39738
rect 10092 39686 10102 39738
rect 10102 39686 10148 39738
rect 9852 39684 9908 39686
rect 9932 39684 9988 39686
rect 10012 39684 10068 39686
rect 10092 39684 10148 39686
rect 9852 38650 9908 38652
rect 9932 38650 9988 38652
rect 10012 38650 10068 38652
rect 10092 38650 10148 38652
rect 9852 38598 9898 38650
rect 9898 38598 9908 38650
rect 9932 38598 9962 38650
rect 9962 38598 9974 38650
rect 9974 38598 9988 38650
rect 10012 38598 10026 38650
rect 10026 38598 10038 38650
rect 10038 38598 10068 38650
rect 10092 38598 10102 38650
rect 10102 38598 10148 38650
rect 9852 38596 9908 38598
rect 9932 38596 9988 38598
rect 10012 38596 10068 38598
rect 10092 38596 10148 38598
rect 9852 37562 9908 37564
rect 9932 37562 9988 37564
rect 10012 37562 10068 37564
rect 10092 37562 10148 37564
rect 9852 37510 9898 37562
rect 9898 37510 9908 37562
rect 9932 37510 9962 37562
rect 9962 37510 9974 37562
rect 9974 37510 9988 37562
rect 10012 37510 10026 37562
rect 10026 37510 10038 37562
rect 10038 37510 10068 37562
rect 10092 37510 10102 37562
rect 10102 37510 10148 37562
rect 9852 37508 9908 37510
rect 9932 37508 9988 37510
rect 10012 37508 10068 37510
rect 10092 37508 10148 37510
rect 9852 36474 9908 36476
rect 9932 36474 9988 36476
rect 10012 36474 10068 36476
rect 10092 36474 10148 36476
rect 9852 36422 9898 36474
rect 9898 36422 9908 36474
rect 9932 36422 9962 36474
rect 9962 36422 9974 36474
rect 9974 36422 9988 36474
rect 10012 36422 10026 36474
rect 10026 36422 10038 36474
rect 10038 36422 10068 36474
rect 10092 36422 10102 36474
rect 10102 36422 10148 36474
rect 9852 36420 9908 36422
rect 9932 36420 9988 36422
rect 10012 36420 10068 36422
rect 10092 36420 10148 36422
rect 9852 35386 9908 35388
rect 9932 35386 9988 35388
rect 10012 35386 10068 35388
rect 10092 35386 10148 35388
rect 9852 35334 9898 35386
rect 9898 35334 9908 35386
rect 9932 35334 9962 35386
rect 9962 35334 9974 35386
rect 9974 35334 9988 35386
rect 10012 35334 10026 35386
rect 10026 35334 10038 35386
rect 10038 35334 10068 35386
rect 10092 35334 10102 35386
rect 10102 35334 10148 35386
rect 9852 35332 9908 35334
rect 9932 35332 9988 35334
rect 10012 35332 10068 35334
rect 10092 35332 10148 35334
rect 9852 34298 9908 34300
rect 9932 34298 9988 34300
rect 10012 34298 10068 34300
rect 10092 34298 10148 34300
rect 9852 34246 9898 34298
rect 9898 34246 9908 34298
rect 9932 34246 9962 34298
rect 9962 34246 9974 34298
rect 9974 34246 9988 34298
rect 10012 34246 10026 34298
rect 10026 34246 10038 34298
rect 10038 34246 10068 34298
rect 10092 34246 10102 34298
rect 10102 34246 10148 34298
rect 9852 34244 9908 34246
rect 9932 34244 9988 34246
rect 10012 34244 10068 34246
rect 10092 34244 10148 34246
rect 9852 33210 9908 33212
rect 9932 33210 9988 33212
rect 10012 33210 10068 33212
rect 10092 33210 10148 33212
rect 9852 33158 9898 33210
rect 9898 33158 9908 33210
rect 9932 33158 9962 33210
rect 9962 33158 9974 33210
rect 9974 33158 9988 33210
rect 10012 33158 10026 33210
rect 10026 33158 10038 33210
rect 10038 33158 10068 33210
rect 10092 33158 10102 33210
rect 10102 33158 10148 33210
rect 9852 33156 9908 33158
rect 9932 33156 9988 33158
rect 10012 33156 10068 33158
rect 10092 33156 10148 33158
rect 12817 44634 12873 44636
rect 12897 44634 12953 44636
rect 12977 44634 13033 44636
rect 13057 44634 13113 44636
rect 12817 44582 12863 44634
rect 12863 44582 12873 44634
rect 12897 44582 12927 44634
rect 12927 44582 12939 44634
rect 12939 44582 12953 44634
rect 12977 44582 12991 44634
rect 12991 44582 13003 44634
rect 13003 44582 13033 44634
rect 13057 44582 13067 44634
rect 13067 44582 13113 44634
rect 12817 44580 12873 44582
rect 12897 44580 12953 44582
rect 12977 44580 13033 44582
rect 13057 44580 13113 44582
rect 15782 45178 15838 45180
rect 15862 45178 15918 45180
rect 15942 45178 15998 45180
rect 16022 45178 16078 45180
rect 15782 45126 15828 45178
rect 15828 45126 15838 45178
rect 15862 45126 15892 45178
rect 15892 45126 15904 45178
rect 15904 45126 15918 45178
rect 15942 45126 15956 45178
rect 15956 45126 15968 45178
rect 15968 45126 15998 45178
rect 16022 45126 16032 45178
rect 16032 45126 16078 45178
rect 15782 45124 15838 45126
rect 15862 45124 15918 45126
rect 15942 45124 15998 45126
rect 16022 45124 16078 45126
rect 9852 32122 9908 32124
rect 9932 32122 9988 32124
rect 10012 32122 10068 32124
rect 10092 32122 10148 32124
rect 9852 32070 9898 32122
rect 9898 32070 9908 32122
rect 9932 32070 9962 32122
rect 9962 32070 9974 32122
rect 9974 32070 9988 32122
rect 10012 32070 10026 32122
rect 10026 32070 10038 32122
rect 10038 32070 10068 32122
rect 10092 32070 10102 32122
rect 10102 32070 10148 32122
rect 9852 32068 9908 32070
rect 9932 32068 9988 32070
rect 10012 32068 10068 32070
rect 10092 32068 10148 32070
rect 9852 31034 9908 31036
rect 9932 31034 9988 31036
rect 10012 31034 10068 31036
rect 10092 31034 10148 31036
rect 9852 30982 9898 31034
rect 9898 30982 9908 31034
rect 9932 30982 9962 31034
rect 9962 30982 9974 31034
rect 9974 30982 9988 31034
rect 10012 30982 10026 31034
rect 10026 30982 10038 31034
rect 10038 30982 10068 31034
rect 10092 30982 10102 31034
rect 10102 30982 10148 31034
rect 9852 30980 9908 30982
rect 9932 30980 9988 30982
rect 10012 30980 10068 30982
rect 10092 30980 10148 30982
rect 9852 29946 9908 29948
rect 9932 29946 9988 29948
rect 10012 29946 10068 29948
rect 10092 29946 10148 29948
rect 9852 29894 9898 29946
rect 9898 29894 9908 29946
rect 9932 29894 9962 29946
rect 9962 29894 9974 29946
rect 9974 29894 9988 29946
rect 10012 29894 10026 29946
rect 10026 29894 10038 29946
rect 10038 29894 10068 29946
rect 10092 29894 10102 29946
rect 10102 29894 10148 29946
rect 9852 29892 9908 29894
rect 9932 29892 9988 29894
rect 10012 29892 10068 29894
rect 10092 29892 10148 29894
rect 9852 28858 9908 28860
rect 9932 28858 9988 28860
rect 10012 28858 10068 28860
rect 10092 28858 10148 28860
rect 9852 28806 9898 28858
rect 9898 28806 9908 28858
rect 9932 28806 9962 28858
rect 9962 28806 9974 28858
rect 9974 28806 9988 28858
rect 10012 28806 10026 28858
rect 10026 28806 10038 28858
rect 10038 28806 10068 28858
rect 10092 28806 10102 28858
rect 10102 28806 10148 28858
rect 9852 28804 9908 28806
rect 9932 28804 9988 28806
rect 10012 28804 10068 28806
rect 10092 28804 10148 28806
rect 9852 27770 9908 27772
rect 9932 27770 9988 27772
rect 10012 27770 10068 27772
rect 10092 27770 10148 27772
rect 9852 27718 9898 27770
rect 9898 27718 9908 27770
rect 9932 27718 9962 27770
rect 9962 27718 9974 27770
rect 9974 27718 9988 27770
rect 10012 27718 10026 27770
rect 10026 27718 10038 27770
rect 10038 27718 10068 27770
rect 10092 27718 10102 27770
rect 10102 27718 10148 27770
rect 9852 27716 9908 27718
rect 9932 27716 9988 27718
rect 10012 27716 10068 27718
rect 10092 27716 10148 27718
rect 9852 26682 9908 26684
rect 9932 26682 9988 26684
rect 10012 26682 10068 26684
rect 10092 26682 10148 26684
rect 9852 26630 9898 26682
rect 9898 26630 9908 26682
rect 9932 26630 9962 26682
rect 9962 26630 9974 26682
rect 9974 26630 9988 26682
rect 10012 26630 10026 26682
rect 10026 26630 10038 26682
rect 10038 26630 10068 26682
rect 10092 26630 10102 26682
rect 10102 26630 10148 26682
rect 9852 26628 9908 26630
rect 9932 26628 9988 26630
rect 10012 26628 10068 26630
rect 10092 26628 10148 26630
rect 9852 25594 9908 25596
rect 9932 25594 9988 25596
rect 10012 25594 10068 25596
rect 10092 25594 10148 25596
rect 9852 25542 9898 25594
rect 9898 25542 9908 25594
rect 9932 25542 9962 25594
rect 9962 25542 9974 25594
rect 9974 25542 9988 25594
rect 10012 25542 10026 25594
rect 10026 25542 10038 25594
rect 10038 25542 10068 25594
rect 10092 25542 10102 25594
rect 10102 25542 10148 25594
rect 9852 25540 9908 25542
rect 9932 25540 9988 25542
rect 10012 25540 10068 25542
rect 10092 25540 10148 25542
rect 9852 24506 9908 24508
rect 9932 24506 9988 24508
rect 10012 24506 10068 24508
rect 10092 24506 10148 24508
rect 9852 24454 9898 24506
rect 9898 24454 9908 24506
rect 9932 24454 9962 24506
rect 9962 24454 9974 24506
rect 9974 24454 9988 24506
rect 10012 24454 10026 24506
rect 10026 24454 10038 24506
rect 10038 24454 10068 24506
rect 10092 24454 10102 24506
rect 10102 24454 10148 24506
rect 9852 24452 9908 24454
rect 9932 24452 9988 24454
rect 10012 24452 10068 24454
rect 10092 24452 10148 24454
rect 9852 23418 9908 23420
rect 9932 23418 9988 23420
rect 10012 23418 10068 23420
rect 10092 23418 10148 23420
rect 9852 23366 9898 23418
rect 9898 23366 9908 23418
rect 9932 23366 9962 23418
rect 9962 23366 9974 23418
rect 9974 23366 9988 23418
rect 10012 23366 10026 23418
rect 10026 23366 10038 23418
rect 10038 23366 10068 23418
rect 10092 23366 10102 23418
rect 10102 23366 10148 23418
rect 9852 23364 9908 23366
rect 9932 23364 9988 23366
rect 10012 23364 10068 23366
rect 10092 23364 10148 23366
rect 6886 17434 6942 17436
rect 6966 17434 7022 17436
rect 7046 17434 7102 17436
rect 7126 17434 7182 17436
rect 6886 17382 6932 17434
rect 6932 17382 6942 17434
rect 6966 17382 6996 17434
rect 6996 17382 7008 17434
rect 7008 17382 7022 17434
rect 7046 17382 7060 17434
rect 7060 17382 7072 17434
rect 7072 17382 7102 17434
rect 7126 17382 7136 17434
rect 7136 17382 7182 17434
rect 6886 17380 6942 17382
rect 6966 17380 7022 17382
rect 7046 17380 7102 17382
rect 7126 17380 7182 17382
rect 6886 16346 6942 16348
rect 6966 16346 7022 16348
rect 7046 16346 7102 16348
rect 7126 16346 7182 16348
rect 6886 16294 6932 16346
rect 6932 16294 6942 16346
rect 6966 16294 6996 16346
rect 6996 16294 7008 16346
rect 7008 16294 7022 16346
rect 7046 16294 7060 16346
rect 7060 16294 7072 16346
rect 7072 16294 7102 16346
rect 7126 16294 7136 16346
rect 7136 16294 7182 16346
rect 6886 16292 6942 16294
rect 6966 16292 7022 16294
rect 7046 16292 7102 16294
rect 7126 16292 7182 16294
rect 7470 15408 7526 15464
rect 3921 8186 3977 8188
rect 4001 8186 4057 8188
rect 4081 8186 4137 8188
rect 4161 8186 4217 8188
rect 3921 8134 3967 8186
rect 3967 8134 3977 8186
rect 4001 8134 4031 8186
rect 4031 8134 4043 8186
rect 4043 8134 4057 8186
rect 4081 8134 4095 8186
rect 4095 8134 4107 8186
rect 4107 8134 4137 8186
rect 4161 8134 4171 8186
rect 4171 8134 4217 8186
rect 3921 8132 3977 8134
rect 4001 8132 4057 8134
rect 4081 8132 4137 8134
rect 4161 8132 4217 8134
rect 3921 7098 3977 7100
rect 4001 7098 4057 7100
rect 4081 7098 4137 7100
rect 4161 7098 4217 7100
rect 3921 7046 3967 7098
rect 3967 7046 3977 7098
rect 4001 7046 4031 7098
rect 4031 7046 4043 7098
rect 4043 7046 4057 7098
rect 4081 7046 4095 7098
rect 4095 7046 4107 7098
rect 4107 7046 4137 7098
rect 4161 7046 4171 7098
rect 4171 7046 4217 7098
rect 3921 7044 3977 7046
rect 4001 7044 4057 7046
rect 4081 7044 4137 7046
rect 4161 7044 4217 7046
rect 3921 6010 3977 6012
rect 4001 6010 4057 6012
rect 4081 6010 4137 6012
rect 4161 6010 4217 6012
rect 3921 5958 3967 6010
rect 3967 5958 3977 6010
rect 4001 5958 4031 6010
rect 4031 5958 4043 6010
rect 4043 5958 4057 6010
rect 4081 5958 4095 6010
rect 4095 5958 4107 6010
rect 4107 5958 4137 6010
rect 4161 5958 4171 6010
rect 4171 5958 4217 6010
rect 3921 5956 3977 5958
rect 4001 5956 4057 5958
rect 4081 5956 4137 5958
rect 4161 5956 4217 5958
rect 3921 4922 3977 4924
rect 4001 4922 4057 4924
rect 4081 4922 4137 4924
rect 4161 4922 4217 4924
rect 3921 4870 3967 4922
rect 3967 4870 3977 4922
rect 4001 4870 4031 4922
rect 4031 4870 4043 4922
rect 4043 4870 4057 4922
rect 4081 4870 4095 4922
rect 4095 4870 4107 4922
rect 4107 4870 4137 4922
rect 4161 4870 4171 4922
rect 4171 4870 4217 4922
rect 3921 4868 3977 4870
rect 4001 4868 4057 4870
rect 4081 4868 4137 4870
rect 4161 4868 4217 4870
rect 6886 15258 6942 15260
rect 6966 15258 7022 15260
rect 7046 15258 7102 15260
rect 7126 15258 7182 15260
rect 6886 15206 6932 15258
rect 6932 15206 6942 15258
rect 6966 15206 6996 15258
rect 6996 15206 7008 15258
rect 7008 15206 7022 15258
rect 7046 15206 7060 15258
rect 7060 15206 7072 15258
rect 7072 15206 7102 15258
rect 7126 15206 7136 15258
rect 7136 15206 7182 15258
rect 6886 15204 6942 15206
rect 6966 15204 7022 15206
rect 7046 15204 7102 15206
rect 7126 15204 7182 15206
rect 6886 14170 6942 14172
rect 6966 14170 7022 14172
rect 7046 14170 7102 14172
rect 7126 14170 7182 14172
rect 6886 14118 6932 14170
rect 6932 14118 6942 14170
rect 6966 14118 6996 14170
rect 6996 14118 7008 14170
rect 7008 14118 7022 14170
rect 7046 14118 7060 14170
rect 7060 14118 7072 14170
rect 7072 14118 7102 14170
rect 7126 14118 7136 14170
rect 7136 14118 7182 14170
rect 6886 14116 6942 14118
rect 6966 14116 7022 14118
rect 7046 14116 7102 14118
rect 7126 14116 7182 14118
rect 6886 13082 6942 13084
rect 6966 13082 7022 13084
rect 7046 13082 7102 13084
rect 7126 13082 7182 13084
rect 6886 13030 6932 13082
rect 6932 13030 6942 13082
rect 6966 13030 6996 13082
rect 6996 13030 7008 13082
rect 7008 13030 7022 13082
rect 7046 13030 7060 13082
rect 7060 13030 7072 13082
rect 7072 13030 7102 13082
rect 7126 13030 7136 13082
rect 7136 13030 7182 13082
rect 6886 13028 6942 13030
rect 6966 13028 7022 13030
rect 7046 13028 7102 13030
rect 7126 13028 7182 13030
rect 6886 11994 6942 11996
rect 6966 11994 7022 11996
rect 7046 11994 7102 11996
rect 7126 11994 7182 11996
rect 6886 11942 6932 11994
rect 6932 11942 6942 11994
rect 6966 11942 6996 11994
rect 6996 11942 7008 11994
rect 7008 11942 7022 11994
rect 7046 11942 7060 11994
rect 7060 11942 7072 11994
rect 7072 11942 7102 11994
rect 7126 11942 7136 11994
rect 7136 11942 7182 11994
rect 6886 11940 6942 11942
rect 6966 11940 7022 11942
rect 7046 11940 7102 11942
rect 7126 11940 7182 11942
rect 9852 22330 9908 22332
rect 9932 22330 9988 22332
rect 10012 22330 10068 22332
rect 10092 22330 10148 22332
rect 9852 22278 9898 22330
rect 9898 22278 9908 22330
rect 9932 22278 9962 22330
rect 9962 22278 9974 22330
rect 9974 22278 9988 22330
rect 10012 22278 10026 22330
rect 10026 22278 10038 22330
rect 10038 22278 10068 22330
rect 10092 22278 10102 22330
rect 10102 22278 10148 22330
rect 9852 22276 9908 22278
rect 9932 22276 9988 22278
rect 10012 22276 10068 22278
rect 10092 22276 10148 22278
rect 12817 43546 12873 43548
rect 12897 43546 12953 43548
rect 12977 43546 13033 43548
rect 13057 43546 13113 43548
rect 12817 43494 12863 43546
rect 12863 43494 12873 43546
rect 12897 43494 12927 43546
rect 12927 43494 12939 43546
rect 12939 43494 12953 43546
rect 12977 43494 12991 43546
rect 12991 43494 13003 43546
rect 13003 43494 13033 43546
rect 13057 43494 13067 43546
rect 13067 43494 13113 43546
rect 12817 43492 12873 43494
rect 12897 43492 12953 43494
rect 12977 43492 13033 43494
rect 13057 43492 13113 43494
rect 12817 42458 12873 42460
rect 12897 42458 12953 42460
rect 12977 42458 13033 42460
rect 13057 42458 13113 42460
rect 12817 42406 12863 42458
rect 12863 42406 12873 42458
rect 12897 42406 12927 42458
rect 12927 42406 12939 42458
rect 12939 42406 12953 42458
rect 12977 42406 12991 42458
rect 12991 42406 13003 42458
rect 13003 42406 13033 42458
rect 13057 42406 13067 42458
rect 13067 42406 13113 42458
rect 12817 42404 12873 42406
rect 12897 42404 12953 42406
rect 12977 42404 13033 42406
rect 13057 42404 13113 42406
rect 12817 41370 12873 41372
rect 12897 41370 12953 41372
rect 12977 41370 13033 41372
rect 13057 41370 13113 41372
rect 12817 41318 12863 41370
rect 12863 41318 12873 41370
rect 12897 41318 12927 41370
rect 12927 41318 12939 41370
rect 12939 41318 12953 41370
rect 12977 41318 12991 41370
rect 12991 41318 13003 41370
rect 13003 41318 13033 41370
rect 13057 41318 13067 41370
rect 13067 41318 13113 41370
rect 12817 41316 12873 41318
rect 12897 41316 12953 41318
rect 12977 41316 13033 41318
rect 13057 41316 13113 41318
rect 12817 40282 12873 40284
rect 12897 40282 12953 40284
rect 12977 40282 13033 40284
rect 13057 40282 13113 40284
rect 12817 40230 12863 40282
rect 12863 40230 12873 40282
rect 12897 40230 12927 40282
rect 12927 40230 12939 40282
rect 12939 40230 12953 40282
rect 12977 40230 12991 40282
rect 12991 40230 13003 40282
rect 13003 40230 13033 40282
rect 13057 40230 13067 40282
rect 13067 40230 13113 40282
rect 12817 40228 12873 40230
rect 12897 40228 12953 40230
rect 12977 40228 13033 40230
rect 13057 40228 13113 40230
rect 12817 39194 12873 39196
rect 12897 39194 12953 39196
rect 12977 39194 13033 39196
rect 13057 39194 13113 39196
rect 12817 39142 12863 39194
rect 12863 39142 12873 39194
rect 12897 39142 12927 39194
rect 12927 39142 12939 39194
rect 12939 39142 12953 39194
rect 12977 39142 12991 39194
rect 12991 39142 13003 39194
rect 13003 39142 13033 39194
rect 13057 39142 13067 39194
rect 13067 39142 13113 39194
rect 12817 39140 12873 39142
rect 12897 39140 12953 39142
rect 12977 39140 13033 39142
rect 13057 39140 13113 39142
rect 12817 38106 12873 38108
rect 12897 38106 12953 38108
rect 12977 38106 13033 38108
rect 13057 38106 13113 38108
rect 12817 38054 12863 38106
rect 12863 38054 12873 38106
rect 12897 38054 12927 38106
rect 12927 38054 12939 38106
rect 12939 38054 12953 38106
rect 12977 38054 12991 38106
rect 12991 38054 13003 38106
rect 13003 38054 13033 38106
rect 13057 38054 13067 38106
rect 13067 38054 13113 38106
rect 12817 38052 12873 38054
rect 12897 38052 12953 38054
rect 12977 38052 13033 38054
rect 13057 38052 13113 38054
rect 15782 44090 15838 44092
rect 15862 44090 15918 44092
rect 15942 44090 15998 44092
rect 16022 44090 16078 44092
rect 15782 44038 15828 44090
rect 15828 44038 15838 44090
rect 15862 44038 15892 44090
rect 15892 44038 15904 44090
rect 15904 44038 15918 44090
rect 15942 44038 15956 44090
rect 15956 44038 15968 44090
rect 15968 44038 15998 44090
rect 16022 44038 16032 44090
rect 16032 44038 16078 44090
rect 15782 44036 15838 44038
rect 15862 44036 15918 44038
rect 15942 44036 15998 44038
rect 16022 44036 16078 44038
rect 15782 43002 15838 43004
rect 15862 43002 15918 43004
rect 15942 43002 15998 43004
rect 16022 43002 16078 43004
rect 15782 42950 15828 43002
rect 15828 42950 15838 43002
rect 15862 42950 15892 43002
rect 15892 42950 15904 43002
rect 15904 42950 15918 43002
rect 15942 42950 15956 43002
rect 15956 42950 15968 43002
rect 15968 42950 15998 43002
rect 16022 42950 16032 43002
rect 16032 42950 16078 43002
rect 15782 42948 15838 42950
rect 15862 42948 15918 42950
rect 15942 42948 15998 42950
rect 16022 42948 16078 42950
rect 15782 41914 15838 41916
rect 15862 41914 15918 41916
rect 15942 41914 15998 41916
rect 16022 41914 16078 41916
rect 15782 41862 15828 41914
rect 15828 41862 15838 41914
rect 15862 41862 15892 41914
rect 15892 41862 15904 41914
rect 15904 41862 15918 41914
rect 15942 41862 15956 41914
rect 15956 41862 15968 41914
rect 15968 41862 15998 41914
rect 16022 41862 16032 41914
rect 16032 41862 16078 41914
rect 15782 41860 15838 41862
rect 15862 41860 15918 41862
rect 15942 41860 15998 41862
rect 16022 41860 16078 41862
rect 12817 37018 12873 37020
rect 12897 37018 12953 37020
rect 12977 37018 13033 37020
rect 13057 37018 13113 37020
rect 12817 36966 12863 37018
rect 12863 36966 12873 37018
rect 12897 36966 12927 37018
rect 12927 36966 12939 37018
rect 12939 36966 12953 37018
rect 12977 36966 12991 37018
rect 12991 36966 13003 37018
rect 13003 36966 13033 37018
rect 13057 36966 13067 37018
rect 13067 36966 13113 37018
rect 12817 36964 12873 36966
rect 12897 36964 12953 36966
rect 12977 36964 13033 36966
rect 13057 36964 13113 36966
rect 12817 35930 12873 35932
rect 12897 35930 12953 35932
rect 12977 35930 13033 35932
rect 13057 35930 13113 35932
rect 12817 35878 12863 35930
rect 12863 35878 12873 35930
rect 12897 35878 12927 35930
rect 12927 35878 12939 35930
rect 12939 35878 12953 35930
rect 12977 35878 12991 35930
rect 12991 35878 13003 35930
rect 13003 35878 13033 35930
rect 13057 35878 13067 35930
rect 13067 35878 13113 35930
rect 12817 35876 12873 35878
rect 12897 35876 12953 35878
rect 12977 35876 13033 35878
rect 13057 35876 13113 35878
rect 12817 34842 12873 34844
rect 12897 34842 12953 34844
rect 12977 34842 13033 34844
rect 13057 34842 13113 34844
rect 12817 34790 12863 34842
rect 12863 34790 12873 34842
rect 12897 34790 12927 34842
rect 12927 34790 12939 34842
rect 12939 34790 12953 34842
rect 12977 34790 12991 34842
rect 12991 34790 13003 34842
rect 13003 34790 13033 34842
rect 13057 34790 13067 34842
rect 13067 34790 13113 34842
rect 12817 34788 12873 34790
rect 12897 34788 12953 34790
rect 12977 34788 13033 34790
rect 13057 34788 13113 34790
rect 12817 33754 12873 33756
rect 12897 33754 12953 33756
rect 12977 33754 13033 33756
rect 13057 33754 13113 33756
rect 12817 33702 12863 33754
rect 12863 33702 12873 33754
rect 12897 33702 12927 33754
rect 12927 33702 12939 33754
rect 12939 33702 12953 33754
rect 12977 33702 12991 33754
rect 12991 33702 13003 33754
rect 13003 33702 13033 33754
rect 13057 33702 13067 33754
rect 13067 33702 13113 33754
rect 12817 33700 12873 33702
rect 12897 33700 12953 33702
rect 12977 33700 13033 33702
rect 13057 33700 13113 33702
rect 12817 32666 12873 32668
rect 12897 32666 12953 32668
rect 12977 32666 13033 32668
rect 13057 32666 13113 32668
rect 12817 32614 12863 32666
rect 12863 32614 12873 32666
rect 12897 32614 12927 32666
rect 12927 32614 12939 32666
rect 12939 32614 12953 32666
rect 12977 32614 12991 32666
rect 12991 32614 13003 32666
rect 13003 32614 13033 32666
rect 13057 32614 13067 32666
rect 13067 32614 13113 32666
rect 12817 32612 12873 32614
rect 12897 32612 12953 32614
rect 12977 32612 13033 32614
rect 13057 32612 13113 32614
rect 9852 21242 9908 21244
rect 9932 21242 9988 21244
rect 10012 21242 10068 21244
rect 10092 21242 10148 21244
rect 9852 21190 9898 21242
rect 9898 21190 9908 21242
rect 9932 21190 9962 21242
rect 9962 21190 9974 21242
rect 9974 21190 9988 21242
rect 10012 21190 10026 21242
rect 10026 21190 10038 21242
rect 10038 21190 10068 21242
rect 10092 21190 10102 21242
rect 10102 21190 10148 21242
rect 9852 21188 9908 21190
rect 9932 21188 9988 21190
rect 10012 21188 10068 21190
rect 10092 21188 10148 21190
rect 6886 10906 6942 10908
rect 6966 10906 7022 10908
rect 7046 10906 7102 10908
rect 7126 10906 7182 10908
rect 6886 10854 6932 10906
rect 6932 10854 6942 10906
rect 6966 10854 6996 10906
rect 6996 10854 7008 10906
rect 7008 10854 7022 10906
rect 7046 10854 7060 10906
rect 7060 10854 7072 10906
rect 7072 10854 7102 10906
rect 7126 10854 7136 10906
rect 7136 10854 7182 10906
rect 6886 10852 6942 10854
rect 6966 10852 7022 10854
rect 7046 10852 7102 10854
rect 7126 10852 7182 10854
rect 7010 10004 7012 10024
rect 7012 10004 7064 10024
rect 7064 10004 7066 10024
rect 7010 9968 7066 10004
rect 6886 9818 6942 9820
rect 6966 9818 7022 9820
rect 7046 9818 7102 9820
rect 7126 9818 7182 9820
rect 6886 9766 6932 9818
rect 6932 9766 6942 9818
rect 6966 9766 6996 9818
rect 6996 9766 7008 9818
rect 7008 9766 7022 9818
rect 7046 9766 7060 9818
rect 7060 9766 7072 9818
rect 7072 9766 7102 9818
rect 7126 9766 7136 9818
rect 7136 9766 7182 9818
rect 6886 9764 6942 9766
rect 6966 9764 7022 9766
rect 7046 9764 7102 9766
rect 7126 9764 7182 9766
rect 7102 9632 7158 9688
rect 6886 8730 6942 8732
rect 6966 8730 7022 8732
rect 7046 8730 7102 8732
rect 7126 8730 7182 8732
rect 6886 8678 6932 8730
rect 6932 8678 6942 8730
rect 6966 8678 6996 8730
rect 6996 8678 7008 8730
rect 7008 8678 7022 8730
rect 7046 8678 7060 8730
rect 7060 8678 7072 8730
rect 7072 8678 7102 8730
rect 7126 8678 7136 8730
rect 7136 8678 7182 8730
rect 6886 8676 6942 8678
rect 6966 8676 7022 8678
rect 7046 8676 7102 8678
rect 7126 8676 7182 8678
rect 6886 7642 6942 7644
rect 6966 7642 7022 7644
rect 7046 7642 7102 7644
rect 7126 7642 7182 7644
rect 6886 7590 6932 7642
rect 6932 7590 6942 7642
rect 6966 7590 6996 7642
rect 6996 7590 7008 7642
rect 7008 7590 7022 7642
rect 7046 7590 7060 7642
rect 7060 7590 7072 7642
rect 7072 7590 7102 7642
rect 7126 7590 7136 7642
rect 7136 7590 7182 7642
rect 6886 7588 6942 7590
rect 6966 7588 7022 7590
rect 7046 7588 7102 7590
rect 7126 7588 7182 7590
rect 6886 6554 6942 6556
rect 6966 6554 7022 6556
rect 7046 6554 7102 6556
rect 7126 6554 7182 6556
rect 6886 6502 6932 6554
rect 6932 6502 6942 6554
rect 6966 6502 6996 6554
rect 6996 6502 7008 6554
rect 7008 6502 7022 6554
rect 7046 6502 7060 6554
rect 7060 6502 7072 6554
rect 7072 6502 7102 6554
rect 7126 6502 7136 6554
rect 7136 6502 7182 6554
rect 6886 6500 6942 6502
rect 6966 6500 7022 6502
rect 7046 6500 7102 6502
rect 7126 6500 7182 6502
rect 6886 5466 6942 5468
rect 6966 5466 7022 5468
rect 7046 5466 7102 5468
rect 7126 5466 7182 5468
rect 6886 5414 6932 5466
rect 6932 5414 6942 5466
rect 6966 5414 6996 5466
rect 6996 5414 7008 5466
rect 7008 5414 7022 5466
rect 7046 5414 7060 5466
rect 7060 5414 7072 5466
rect 7072 5414 7102 5466
rect 7126 5414 7136 5466
rect 7136 5414 7182 5466
rect 6886 5412 6942 5414
rect 6966 5412 7022 5414
rect 7046 5412 7102 5414
rect 7126 5412 7182 5414
rect 9852 20154 9908 20156
rect 9932 20154 9988 20156
rect 10012 20154 10068 20156
rect 10092 20154 10148 20156
rect 9852 20102 9898 20154
rect 9898 20102 9908 20154
rect 9932 20102 9962 20154
rect 9962 20102 9974 20154
rect 9974 20102 9988 20154
rect 10012 20102 10026 20154
rect 10026 20102 10038 20154
rect 10038 20102 10068 20154
rect 10092 20102 10102 20154
rect 10102 20102 10148 20154
rect 9852 20100 9908 20102
rect 9932 20100 9988 20102
rect 10012 20100 10068 20102
rect 10092 20100 10148 20102
rect 9852 19066 9908 19068
rect 9932 19066 9988 19068
rect 10012 19066 10068 19068
rect 10092 19066 10148 19068
rect 9852 19014 9898 19066
rect 9898 19014 9908 19066
rect 9932 19014 9962 19066
rect 9962 19014 9974 19066
rect 9974 19014 9988 19066
rect 10012 19014 10026 19066
rect 10026 19014 10038 19066
rect 10038 19014 10068 19066
rect 10092 19014 10102 19066
rect 10102 19014 10148 19066
rect 9852 19012 9908 19014
rect 9932 19012 9988 19014
rect 10012 19012 10068 19014
rect 10092 19012 10148 19014
rect 9852 17978 9908 17980
rect 9932 17978 9988 17980
rect 10012 17978 10068 17980
rect 10092 17978 10148 17980
rect 9852 17926 9898 17978
rect 9898 17926 9908 17978
rect 9932 17926 9962 17978
rect 9962 17926 9974 17978
rect 9974 17926 9988 17978
rect 10012 17926 10026 17978
rect 10026 17926 10038 17978
rect 10038 17926 10068 17978
rect 10092 17926 10102 17978
rect 10102 17926 10148 17978
rect 9852 17924 9908 17926
rect 9932 17924 9988 17926
rect 10012 17924 10068 17926
rect 10092 17924 10148 17926
rect 9852 16890 9908 16892
rect 9932 16890 9988 16892
rect 10012 16890 10068 16892
rect 10092 16890 10148 16892
rect 9852 16838 9898 16890
rect 9898 16838 9908 16890
rect 9932 16838 9962 16890
rect 9962 16838 9974 16890
rect 9974 16838 9988 16890
rect 10012 16838 10026 16890
rect 10026 16838 10038 16890
rect 10038 16838 10068 16890
rect 10092 16838 10102 16890
rect 10102 16838 10148 16890
rect 9852 16836 9908 16838
rect 9932 16836 9988 16838
rect 10012 16836 10068 16838
rect 10092 16836 10148 16838
rect 9852 15802 9908 15804
rect 9932 15802 9988 15804
rect 10012 15802 10068 15804
rect 10092 15802 10148 15804
rect 9852 15750 9898 15802
rect 9898 15750 9908 15802
rect 9932 15750 9962 15802
rect 9962 15750 9974 15802
rect 9974 15750 9988 15802
rect 10012 15750 10026 15802
rect 10026 15750 10038 15802
rect 10038 15750 10068 15802
rect 10092 15750 10102 15802
rect 10102 15750 10148 15802
rect 9852 15748 9908 15750
rect 9932 15748 9988 15750
rect 10012 15748 10068 15750
rect 10092 15748 10148 15750
rect 9852 14714 9908 14716
rect 9932 14714 9988 14716
rect 10012 14714 10068 14716
rect 10092 14714 10148 14716
rect 9852 14662 9898 14714
rect 9898 14662 9908 14714
rect 9932 14662 9962 14714
rect 9962 14662 9974 14714
rect 9974 14662 9988 14714
rect 10012 14662 10026 14714
rect 10026 14662 10038 14714
rect 10038 14662 10068 14714
rect 10092 14662 10102 14714
rect 10102 14662 10148 14714
rect 9852 14660 9908 14662
rect 9932 14660 9988 14662
rect 10012 14660 10068 14662
rect 10092 14660 10148 14662
rect 9852 13626 9908 13628
rect 9932 13626 9988 13628
rect 10012 13626 10068 13628
rect 10092 13626 10148 13628
rect 9852 13574 9898 13626
rect 9898 13574 9908 13626
rect 9932 13574 9962 13626
rect 9962 13574 9974 13626
rect 9974 13574 9988 13626
rect 10012 13574 10026 13626
rect 10026 13574 10038 13626
rect 10038 13574 10068 13626
rect 10092 13574 10102 13626
rect 10102 13574 10148 13626
rect 9852 13572 9908 13574
rect 9932 13572 9988 13574
rect 10012 13572 10068 13574
rect 10092 13572 10148 13574
rect 9852 12538 9908 12540
rect 9932 12538 9988 12540
rect 10012 12538 10068 12540
rect 10092 12538 10148 12540
rect 9852 12486 9898 12538
rect 9898 12486 9908 12538
rect 9932 12486 9962 12538
rect 9962 12486 9974 12538
rect 9974 12486 9988 12538
rect 10012 12486 10026 12538
rect 10026 12486 10038 12538
rect 10038 12486 10068 12538
rect 10092 12486 10102 12538
rect 10102 12486 10148 12538
rect 9852 12484 9908 12486
rect 9932 12484 9988 12486
rect 10012 12484 10068 12486
rect 10092 12484 10148 12486
rect 3921 3834 3977 3836
rect 4001 3834 4057 3836
rect 4081 3834 4137 3836
rect 4161 3834 4217 3836
rect 3921 3782 3967 3834
rect 3967 3782 3977 3834
rect 4001 3782 4031 3834
rect 4031 3782 4043 3834
rect 4043 3782 4057 3834
rect 4081 3782 4095 3834
rect 4095 3782 4107 3834
rect 4107 3782 4137 3834
rect 4161 3782 4171 3834
rect 4171 3782 4217 3834
rect 3921 3780 3977 3782
rect 4001 3780 4057 3782
rect 4081 3780 4137 3782
rect 4161 3780 4217 3782
rect 6886 4378 6942 4380
rect 6966 4378 7022 4380
rect 7046 4378 7102 4380
rect 7126 4378 7182 4380
rect 6886 4326 6932 4378
rect 6932 4326 6942 4378
rect 6966 4326 6996 4378
rect 6996 4326 7008 4378
rect 7008 4326 7022 4378
rect 7046 4326 7060 4378
rect 7060 4326 7072 4378
rect 7072 4326 7102 4378
rect 7126 4326 7136 4378
rect 7136 4326 7182 4378
rect 6886 4324 6942 4326
rect 6966 4324 7022 4326
rect 7046 4324 7102 4326
rect 7126 4324 7182 4326
rect 8758 9968 8814 10024
rect 9852 11450 9908 11452
rect 9932 11450 9988 11452
rect 10012 11450 10068 11452
rect 10092 11450 10148 11452
rect 9852 11398 9898 11450
rect 9898 11398 9908 11450
rect 9932 11398 9962 11450
rect 9962 11398 9974 11450
rect 9974 11398 9988 11450
rect 10012 11398 10026 11450
rect 10026 11398 10038 11450
rect 10038 11398 10068 11450
rect 10092 11398 10102 11450
rect 10102 11398 10148 11450
rect 9852 11396 9908 11398
rect 9932 11396 9988 11398
rect 10012 11396 10068 11398
rect 10092 11396 10148 11398
rect 12817 31578 12873 31580
rect 12897 31578 12953 31580
rect 12977 31578 13033 31580
rect 13057 31578 13113 31580
rect 12817 31526 12863 31578
rect 12863 31526 12873 31578
rect 12897 31526 12927 31578
rect 12927 31526 12939 31578
rect 12939 31526 12953 31578
rect 12977 31526 12991 31578
rect 12991 31526 13003 31578
rect 13003 31526 13033 31578
rect 13057 31526 13067 31578
rect 13067 31526 13113 31578
rect 12817 31524 12873 31526
rect 12897 31524 12953 31526
rect 12977 31524 13033 31526
rect 13057 31524 13113 31526
rect 12817 30490 12873 30492
rect 12897 30490 12953 30492
rect 12977 30490 13033 30492
rect 13057 30490 13113 30492
rect 12817 30438 12863 30490
rect 12863 30438 12873 30490
rect 12897 30438 12927 30490
rect 12927 30438 12939 30490
rect 12939 30438 12953 30490
rect 12977 30438 12991 30490
rect 12991 30438 13003 30490
rect 13003 30438 13033 30490
rect 13057 30438 13067 30490
rect 13067 30438 13113 30490
rect 12817 30436 12873 30438
rect 12897 30436 12953 30438
rect 12977 30436 13033 30438
rect 13057 30436 13113 30438
rect 12817 29402 12873 29404
rect 12897 29402 12953 29404
rect 12977 29402 13033 29404
rect 13057 29402 13113 29404
rect 12817 29350 12863 29402
rect 12863 29350 12873 29402
rect 12897 29350 12927 29402
rect 12927 29350 12939 29402
rect 12939 29350 12953 29402
rect 12977 29350 12991 29402
rect 12991 29350 13003 29402
rect 13003 29350 13033 29402
rect 13057 29350 13067 29402
rect 13067 29350 13113 29402
rect 12817 29348 12873 29350
rect 12897 29348 12953 29350
rect 12977 29348 13033 29350
rect 13057 29348 13113 29350
rect 9852 10362 9908 10364
rect 9932 10362 9988 10364
rect 10012 10362 10068 10364
rect 10092 10362 10148 10364
rect 9852 10310 9898 10362
rect 9898 10310 9908 10362
rect 9932 10310 9962 10362
rect 9962 10310 9974 10362
rect 9974 10310 9988 10362
rect 10012 10310 10026 10362
rect 10026 10310 10038 10362
rect 10038 10310 10068 10362
rect 10092 10310 10102 10362
rect 10102 10310 10148 10362
rect 9852 10308 9908 10310
rect 9932 10308 9988 10310
rect 10012 10308 10068 10310
rect 10092 10308 10148 10310
rect 9852 9274 9908 9276
rect 9932 9274 9988 9276
rect 10012 9274 10068 9276
rect 10092 9274 10148 9276
rect 9852 9222 9898 9274
rect 9898 9222 9908 9274
rect 9932 9222 9962 9274
rect 9962 9222 9974 9274
rect 9974 9222 9988 9274
rect 10012 9222 10026 9274
rect 10026 9222 10038 9274
rect 10038 9222 10068 9274
rect 10092 9222 10102 9274
rect 10102 9222 10148 9274
rect 9852 9220 9908 9222
rect 9932 9220 9988 9222
rect 10012 9220 10068 9222
rect 10092 9220 10148 9222
rect 9852 8186 9908 8188
rect 9932 8186 9988 8188
rect 10012 8186 10068 8188
rect 10092 8186 10148 8188
rect 9852 8134 9898 8186
rect 9898 8134 9908 8186
rect 9932 8134 9962 8186
rect 9962 8134 9974 8186
rect 9974 8134 9988 8186
rect 10012 8134 10026 8186
rect 10026 8134 10038 8186
rect 10038 8134 10068 8186
rect 10092 8134 10102 8186
rect 10102 8134 10148 8186
rect 9852 8132 9908 8134
rect 9932 8132 9988 8134
rect 10012 8132 10068 8134
rect 10092 8132 10148 8134
rect 9852 7098 9908 7100
rect 9932 7098 9988 7100
rect 10012 7098 10068 7100
rect 10092 7098 10148 7100
rect 9852 7046 9898 7098
rect 9898 7046 9908 7098
rect 9932 7046 9962 7098
rect 9962 7046 9974 7098
rect 9974 7046 9988 7098
rect 10012 7046 10026 7098
rect 10026 7046 10038 7098
rect 10038 7046 10068 7098
rect 10092 7046 10102 7098
rect 10102 7046 10148 7098
rect 9852 7044 9908 7046
rect 9932 7044 9988 7046
rect 10012 7044 10068 7046
rect 10092 7044 10148 7046
rect 9852 6010 9908 6012
rect 9932 6010 9988 6012
rect 10012 6010 10068 6012
rect 10092 6010 10148 6012
rect 9852 5958 9898 6010
rect 9898 5958 9908 6010
rect 9932 5958 9962 6010
rect 9962 5958 9974 6010
rect 9974 5958 9988 6010
rect 10012 5958 10026 6010
rect 10026 5958 10038 6010
rect 10038 5958 10068 6010
rect 10092 5958 10102 6010
rect 10102 5958 10148 6010
rect 9852 5956 9908 5958
rect 9932 5956 9988 5958
rect 10012 5956 10068 5958
rect 10092 5956 10148 5958
rect 9852 4922 9908 4924
rect 9932 4922 9988 4924
rect 10012 4922 10068 4924
rect 10092 4922 10148 4924
rect 9852 4870 9898 4922
rect 9898 4870 9908 4922
rect 9932 4870 9962 4922
rect 9962 4870 9974 4922
rect 9974 4870 9988 4922
rect 10012 4870 10026 4922
rect 10026 4870 10038 4922
rect 10038 4870 10068 4922
rect 10092 4870 10102 4922
rect 10102 4870 10148 4922
rect 9852 4868 9908 4870
rect 9932 4868 9988 4870
rect 10012 4868 10068 4870
rect 10092 4868 10148 4870
rect 9852 3834 9908 3836
rect 9932 3834 9988 3836
rect 10012 3834 10068 3836
rect 10092 3834 10148 3836
rect 9852 3782 9898 3834
rect 9898 3782 9908 3834
rect 9932 3782 9962 3834
rect 9962 3782 9974 3834
rect 9974 3782 9988 3834
rect 10012 3782 10026 3834
rect 10026 3782 10038 3834
rect 10038 3782 10068 3834
rect 10092 3782 10102 3834
rect 10102 3782 10148 3834
rect 9852 3780 9908 3782
rect 9932 3780 9988 3782
rect 10012 3780 10068 3782
rect 10092 3780 10148 3782
rect 12817 28314 12873 28316
rect 12897 28314 12953 28316
rect 12977 28314 13033 28316
rect 13057 28314 13113 28316
rect 12817 28262 12863 28314
rect 12863 28262 12873 28314
rect 12897 28262 12927 28314
rect 12927 28262 12939 28314
rect 12939 28262 12953 28314
rect 12977 28262 12991 28314
rect 12991 28262 13003 28314
rect 13003 28262 13033 28314
rect 13057 28262 13067 28314
rect 13067 28262 13113 28314
rect 12817 28260 12873 28262
rect 12897 28260 12953 28262
rect 12977 28260 13033 28262
rect 13057 28260 13113 28262
rect 12817 27226 12873 27228
rect 12897 27226 12953 27228
rect 12977 27226 13033 27228
rect 13057 27226 13113 27228
rect 12817 27174 12863 27226
rect 12863 27174 12873 27226
rect 12897 27174 12927 27226
rect 12927 27174 12939 27226
rect 12939 27174 12953 27226
rect 12977 27174 12991 27226
rect 12991 27174 13003 27226
rect 13003 27174 13033 27226
rect 13057 27174 13067 27226
rect 13067 27174 13113 27226
rect 12817 27172 12873 27174
rect 12897 27172 12953 27174
rect 12977 27172 13033 27174
rect 13057 27172 13113 27174
rect 15782 40826 15838 40828
rect 15862 40826 15918 40828
rect 15942 40826 15998 40828
rect 16022 40826 16078 40828
rect 15782 40774 15828 40826
rect 15828 40774 15838 40826
rect 15862 40774 15892 40826
rect 15892 40774 15904 40826
rect 15904 40774 15918 40826
rect 15942 40774 15956 40826
rect 15956 40774 15968 40826
rect 15968 40774 15998 40826
rect 16022 40774 16032 40826
rect 16032 40774 16078 40826
rect 15782 40772 15838 40774
rect 15862 40772 15918 40774
rect 15942 40772 15998 40774
rect 16022 40772 16078 40774
rect 15782 39738 15838 39740
rect 15862 39738 15918 39740
rect 15942 39738 15998 39740
rect 16022 39738 16078 39740
rect 15782 39686 15828 39738
rect 15828 39686 15838 39738
rect 15862 39686 15892 39738
rect 15892 39686 15904 39738
rect 15904 39686 15918 39738
rect 15942 39686 15956 39738
rect 15956 39686 15968 39738
rect 15968 39686 15998 39738
rect 16022 39686 16032 39738
rect 16032 39686 16078 39738
rect 15782 39684 15838 39686
rect 15862 39684 15918 39686
rect 15942 39684 15998 39686
rect 16022 39684 16078 39686
rect 15782 38650 15838 38652
rect 15862 38650 15918 38652
rect 15942 38650 15998 38652
rect 16022 38650 16078 38652
rect 15782 38598 15828 38650
rect 15828 38598 15838 38650
rect 15862 38598 15892 38650
rect 15892 38598 15904 38650
rect 15904 38598 15918 38650
rect 15942 38598 15956 38650
rect 15956 38598 15968 38650
rect 15968 38598 15998 38650
rect 16022 38598 16032 38650
rect 16032 38598 16078 38650
rect 15782 38596 15838 38598
rect 15862 38596 15918 38598
rect 15942 38596 15998 38598
rect 16022 38596 16078 38598
rect 15782 37562 15838 37564
rect 15862 37562 15918 37564
rect 15942 37562 15998 37564
rect 16022 37562 16078 37564
rect 15782 37510 15828 37562
rect 15828 37510 15838 37562
rect 15862 37510 15892 37562
rect 15892 37510 15904 37562
rect 15904 37510 15918 37562
rect 15942 37510 15956 37562
rect 15956 37510 15968 37562
rect 15968 37510 15998 37562
rect 16022 37510 16032 37562
rect 16032 37510 16078 37562
rect 15782 37508 15838 37510
rect 15862 37508 15918 37510
rect 15942 37508 15998 37510
rect 16022 37508 16078 37510
rect 15782 36474 15838 36476
rect 15862 36474 15918 36476
rect 15942 36474 15998 36476
rect 16022 36474 16078 36476
rect 15782 36422 15828 36474
rect 15828 36422 15838 36474
rect 15862 36422 15892 36474
rect 15892 36422 15904 36474
rect 15904 36422 15918 36474
rect 15942 36422 15956 36474
rect 15956 36422 15968 36474
rect 15968 36422 15998 36474
rect 16022 36422 16032 36474
rect 16032 36422 16078 36474
rect 15782 36420 15838 36422
rect 15862 36420 15918 36422
rect 15942 36420 15998 36422
rect 16022 36420 16078 36422
rect 18142 40840 18198 40896
rect 15782 35386 15838 35388
rect 15862 35386 15918 35388
rect 15942 35386 15998 35388
rect 16022 35386 16078 35388
rect 15782 35334 15828 35386
rect 15828 35334 15838 35386
rect 15862 35334 15892 35386
rect 15892 35334 15904 35386
rect 15904 35334 15918 35386
rect 15942 35334 15956 35386
rect 15956 35334 15968 35386
rect 15968 35334 15998 35386
rect 16022 35334 16032 35386
rect 16032 35334 16078 35386
rect 15782 35332 15838 35334
rect 15862 35332 15918 35334
rect 15942 35332 15998 35334
rect 16022 35332 16078 35334
rect 15782 34298 15838 34300
rect 15862 34298 15918 34300
rect 15942 34298 15998 34300
rect 16022 34298 16078 34300
rect 15782 34246 15828 34298
rect 15828 34246 15838 34298
rect 15862 34246 15892 34298
rect 15892 34246 15904 34298
rect 15904 34246 15918 34298
rect 15942 34246 15956 34298
rect 15956 34246 15968 34298
rect 15968 34246 15998 34298
rect 16022 34246 16032 34298
rect 16032 34246 16078 34298
rect 15782 34244 15838 34246
rect 15862 34244 15918 34246
rect 15942 34244 15998 34246
rect 16022 34244 16078 34246
rect 15782 33210 15838 33212
rect 15862 33210 15918 33212
rect 15942 33210 15998 33212
rect 16022 33210 16078 33212
rect 15782 33158 15828 33210
rect 15828 33158 15838 33210
rect 15862 33158 15892 33210
rect 15892 33158 15904 33210
rect 15904 33158 15918 33210
rect 15942 33158 15956 33210
rect 15956 33158 15968 33210
rect 15968 33158 15998 33210
rect 16022 33158 16032 33210
rect 16032 33158 16078 33210
rect 15782 33156 15838 33158
rect 15862 33156 15918 33158
rect 15942 33156 15998 33158
rect 16022 33156 16078 33158
rect 12817 26138 12873 26140
rect 12897 26138 12953 26140
rect 12977 26138 13033 26140
rect 13057 26138 13113 26140
rect 12817 26086 12863 26138
rect 12863 26086 12873 26138
rect 12897 26086 12927 26138
rect 12927 26086 12939 26138
rect 12939 26086 12953 26138
rect 12977 26086 12991 26138
rect 12991 26086 13003 26138
rect 13003 26086 13033 26138
rect 13057 26086 13067 26138
rect 13067 26086 13113 26138
rect 12817 26084 12873 26086
rect 12897 26084 12953 26086
rect 12977 26084 13033 26086
rect 13057 26084 13113 26086
rect 12817 25050 12873 25052
rect 12897 25050 12953 25052
rect 12977 25050 13033 25052
rect 13057 25050 13113 25052
rect 12817 24998 12863 25050
rect 12863 24998 12873 25050
rect 12897 24998 12927 25050
rect 12927 24998 12939 25050
rect 12939 24998 12953 25050
rect 12977 24998 12991 25050
rect 12991 24998 13003 25050
rect 13003 24998 13033 25050
rect 13057 24998 13067 25050
rect 13067 24998 13113 25050
rect 12817 24996 12873 24998
rect 12897 24996 12953 24998
rect 12977 24996 13033 24998
rect 13057 24996 13113 24998
rect 12817 23962 12873 23964
rect 12897 23962 12953 23964
rect 12977 23962 13033 23964
rect 13057 23962 13113 23964
rect 12817 23910 12863 23962
rect 12863 23910 12873 23962
rect 12897 23910 12927 23962
rect 12927 23910 12939 23962
rect 12939 23910 12953 23962
rect 12977 23910 12991 23962
rect 12991 23910 13003 23962
rect 13003 23910 13033 23962
rect 13057 23910 13067 23962
rect 13067 23910 13113 23962
rect 12817 23908 12873 23910
rect 12897 23908 12953 23910
rect 12977 23908 13033 23910
rect 13057 23908 13113 23910
rect 12817 22874 12873 22876
rect 12897 22874 12953 22876
rect 12977 22874 13033 22876
rect 13057 22874 13113 22876
rect 12817 22822 12863 22874
rect 12863 22822 12873 22874
rect 12897 22822 12927 22874
rect 12927 22822 12939 22874
rect 12939 22822 12953 22874
rect 12977 22822 12991 22874
rect 12991 22822 13003 22874
rect 13003 22822 13033 22874
rect 13057 22822 13067 22874
rect 13067 22822 13113 22874
rect 12817 22820 12873 22822
rect 12897 22820 12953 22822
rect 12977 22820 13033 22822
rect 13057 22820 13113 22822
rect 12817 21786 12873 21788
rect 12897 21786 12953 21788
rect 12977 21786 13033 21788
rect 13057 21786 13113 21788
rect 12817 21734 12863 21786
rect 12863 21734 12873 21786
rect 12897 21734 12927 21786
rect 12927 21734 12939 21786
rect 12939 21734 12953 21786
rect 12977 21734 12991 21786
rect 12991 21734 13003 21786
rect 13003 21734 13033 21786
rect 13057 21734 13067 21786
rect 13067 21734 13113 21786
rect 12817 21732 12873 21734
rect 12897 21732 12953 21734
rect 12977 21732 13033 21734
rect 13057 21732 13113 21734
rect 12817 20698 12873 20700
rect 12897 20698 12953 20700
rect 12977 20698 13033 20700
rect 13057 20698 13113 20700
rect 12817 20646 12863 20698
rect 12863 20646 12873 20698
rect 12897 20646 12927 20698
rect 12927 20646 12939 20698
rect 12939 20646 12953 20698
rect 12977 20646 12991 20698
rect 12991 20646 13003 20698
rect 13003 20646 13033 20698
rect 13057 20646 13067 20698
rect 13067 20646 13113 20698
rect 12817 20644 12873 20646
rect 12897 20644 12953 20646
rect 12977 20644 13033 20646
rect 13057 20644 13113 20646
rect 12817 19610 12873 19612
rect 12897 19610 12953 19612
rect 12977 19610 13033 19612
rect 13057 19610 13113 19612
rect 12817 19558 12863 19610
rect 12863 19558 12873 19610
rect 12897 19558 12927 19610
rect 12927 19558 12939 19610
rect 12939 19558 12953 19610
rect 12977 19558 12991 19610
rect 12991 19558 13003 19610
rect 13003 19558 13033 19610
rect 13057 19558 13067 19610
rect 13067 19558 13113 19610
rect 12817 19556 12873 19558
rect 12897 19556 12953 19558
rect 12977 19556 13033 19558
rect 13057 19556 13113 19558
rect 12817 18522 12873 18524
rect 12897 18522 12953 18524
rect 12977 18522 13033 18524
rect 13057 18522 13113 18524
rect 12817 18470 12863 18522
rect 12863 18470 12873 18522
rect 12897 18470 12927 18522
rect 12927 18470 12939 18522
rect 12939 18470 12953 18522
rect 12977 18470 12991 18522
rect 12991 18470 13003 18522
rect 13003 18470 13033 18522
rect 13057 18470 13067 18522
rect 13067 18470 13113 18522
rect 12817 18468 12873 18470
rect 12897 18468 12953 18470
rect 12977 18468 13033 18470
rect 13057 18468 13113 18470
rect 12817 17434 12873 17436
rect 12897 17434 12953 17436
rect 12977 17434 13033 17436
rect 13057 17434 13113 17436
rect 12817 17382 12863 17434
rect 12863 17382 12873 17434
rect 12897 17382 12927 17434
rect 12927 17382 12939 17434
rect 12939 17382 12953 17434
rect 12977 17382 12991 17434
rect 12991 17382 13003 17434
rect 13003 17382 13033 17434
rect 13057 17382 13067 17434
rect 13067 17382 13113 17434
rect 12817 17380 12873 17382
rect 12897 17380 12953 17382
rect 12977 17380 13033 17382
rect 13057 17380 13113 17382
rect 12817 16346 12873 16348
rect 12897 16346 12953 16348
rect 12977 16346 13033 16348
rect 13057 16346 13113 16348
rect 12817 16294 12863 16346
rect 12863 16294 12873 16346
rect 12897 16294 12927 16346
rect 12927 16294 12939 16346
rect 12939 16294 12953 16346
rect 12977 16294 12991 16346
rect 12991 16294 13003 16346
rect 13003 16294 13033 16346
rect 13057 16294 13067 16346
rect 13067 16294 13113 16346
rect 12817 16292 12873 16294
rect 12897 16292 12953 16294
rect 12977 16292 13033 16294
rect 13057 16292 13113 16294
rect 12817 15258 12873 15260
rect 12897 15258 12953 15260
rect 12977 15258 13033 15260
rect 13057 15258 13113 15260
rect 12817 15206 12863 15258
rect 12863 15206 12873 15258
rect 12897 15206 12927 15258
rect 12927 15206 12939 15258
rect 12939 15206 12953 15258
rect 12977 15206 12991 15258
rect 12991 15206 13003 15258
rect 13003 15206 13033 15258
rect 13057 15206 13067 15258
rect 13067 15206 13113 15258
rect 12817 15204 12873 15206
rect 12897 15204 12953 15206
rect 12977 15204 13033 15206
rect 13057 15204 13113 15206
rect 12817 14170 12873 14172
rect 12897 14170 12953 14172
rect 12977 14170 13033 14172
rect 13057 14170 13113 14172
rect 12817 14118 12863 14170
rect 12863 14118 12873 14170
rect 12897 14118 12927 14170
rect 12927 14118 12939 14170
rect 12939 14118 12953 14170
rect 12977 14118 12991 14170
rect 12991 14118 13003 14170
rect 13003 14118 13033 14170
rect 13057 14118 13067 14170
rect 13067 14118 13113 14170
rect 12817 14116 12873 14118
rect 12897 14116 12953 14118
rect 12977 14116 13033 14118
rect 13057 14116 13113 14118
rect 12817 13082 12873 13084
rect 12897 13082 12953 13084
rect 12977 13082 13033 13084
rect 13057 13082 13113 13084
rect 12817 13030 12863 13082
rect 12863 13030 12873 13082
rect 12897 13030 12927 13082
rect 12927 13030 12939 13082
rect 12939 13030 12953 13082
rect 12977 13030 12991 13082
rect 12991 13030 13003 13082
rect 13003 13030 13033 13082
rect 13057 13030 13067 13082
rect 13067 13030 13113 13082
rect 12817 13028 12873 13030
rect 12897 13028 12953 13030
rect 12977 13028 13033 13030
rect 13057 13028 13113 13030
rect 15782 32122 15838 32124
rect 15862 32122 15918 32124
rect 15942 32122 15998 32124
rect 16022 32122 16078 32124
rect 15782 32070 15828 32122
rect 15828 32070 15838 32122
rect 15862 32070 15892 32122
rect 15892 32070 15904 32122
rect 15904 32070 15918 32122
rect 15942 32070 15956 32122
rect 15956 32070 15968 32122
rect 15968 32070 15998 32122
rect 16022 32070 16032 32122
rect 16032 32070 16078 32122
rect 15782 32068 15838 32070
rect 15862 32068 15918 32070
rect 15942 32068 15998 32070
rect 16022 32068 16078 32070
rect 15782 31034 15838 31036
rect 15862 31034 15918 31036
rect 15942 31034 15998 31036
rect 16022 31034 16078 31036
rect 15782 30982 15828 31034
rect 15828 30982 15838 31034
rect 15862 30982 15892 31034
rect 15892 30982 15904 31034
rect 15904 30982 15918 31034
rect 15942 30982 15956 31034
rect 15956 30982 15968 31034
rect 15968 30982 15998 31034
rect 16022 30982 16032 31034
rect 16032 30982 16078 31034
rect 15782 30980 15838 30982
rect 15862 30980 15918 30982
rect 15942 30980 15998 30982
rect 16022 30980 16078 30982
rect 15782 29946 15838 29948
rect 15862 29946 15918 29948
rect 15942 29946 15998 29948
rect 16022 29946 16078 29948
rect 15782 29894 15828 29946
rect 15828 29894 15838 29946
rect 15862 29894 15892 29946
rect 15892 29894 15904 29946
rect 15904 29894 15918 29946
rect 15942 29894 15956 29946
rect 15956 29894 15968 29946
rect 15968 29894 15998 29946
rect 16022 29894 16032 29946
rect 16032 29894 16078 29946
rect 15782 29892 15838 29894
rect 15862 29892 15918 29894
rect 15942 29892 15998 29894
rect 16022 29892 16078 29894
rect 15782 28858 15838 28860
rect 15862 28858 15918 28860
rect 15942 28858 15998 28860
rect 16022 28858 16078 28860
rect 15782 28806 15828 28858
rect 15828 28806 15838 28858
rect 15862 28806 15892 28858
rect 15892 28806 15904 28858
rect 15904 28806 15918 28858
rect 15942 28806 15956 28858
rect 15956 28806 15968 28858
rect 15968 28806 15998 28858
rect 16022 28806 16032 28858
rect 16032 28806 16078 28858
rect 15782 28804 15838 28806
rect 15862 28804 15918 28806
rect 15942 28804 15998 28806
rect 16022 28804 16078 28806
rect 15782 27770 15838 27772
rect 15862 27770 15918 27772
rect 15942 27770 15998 27772
rect 16022 27770 16078 27772
rect 15782 27718 15828 27770
rect 15828 27718 15838 27770
rect 15862 27718 15892 27770
rect 15892 27718 15904 27770
rect 15904 27718 15918 27770
rect 15942 27718 15956 27770
rect 15956 27718 15968 27770
rect 15968 27718 15998 27770
rect 16022 27718 16032 27770
rect 16032 27718 16078 27770
rect 15782 27716 15838 27718
rect 15862 27716 15918 27718
rect 15942 27716 15998 27718
rect 16022 27716 16078 27718
rect 15782 26682 15838 26684
rect 15862 26682 15918 26684
rect 15942 26682 15998 26684
rect 16022 26682 16078 26684
rect 15782 26630 15828 26682
rect 15828 26630 15838 26682
rect 15862 26630 15892 26682
rect 15892 26630 15904 26682
rect 15904 26630 15918 26682
rect 15942 26630 15956 26682
rect 15956 26630 15968 26682
rect 15968 26630 15998 26682
rect 16022 26630 16032 26682
rect 16032 26630 16078 26682
rect 15782 26628 15838 26630
rect 15862 26628 15918 26630
rect 15942 26628 15998 26630
rect 16022 26628 16078 26630
rect 15782 25594 15838 25596
rect 15862 25594 15918 25596
rect 15942 25594 15998 25596
rect 16022 25594 16078 25596
rect 15782 25542 15828 25594
rect 15828 25542 15838 25594
rect 15862 25542 15892 25594
rect 15892 25542 15904 25594
rect 15904 25542 15918 25594
rect 15942 25542 15956 25594
rect 15956 25542 15968 25594
rect 15968 25542 15998 25594
rect 16022 25542 16032 25594
rect 16032 25542 16078 25594
rect 15782 25540 15838 25542
rect 15862 25540 15918 25542
rect 15942 25540 15998 25542
rect 16022 25540 16078 25542
rect 15782 24506 15838 24508
rect 15862 24506 15918 24508
rect 15942 24506 15998 24508
rect 16022 24506 16078 24508
rect 15782 24454 15828 24506
rect 15828 24454 15838 24506
rect 15862 24454 15892 24506
rect 15892 24454 15904 24506
rect 15904 24454 15918 24506
rect 15942 24454 15956 24506
rect 15956 24454 15968 24506
rect 15968 24454 15998 24506
rect 16022 24454 16032 24506
rect 16032 24454 16078 24506
rect 15782 24452 15838 24454
rect 15862 24452 15918 24454
rect 15942 24452 15998 24454
rect 16022 24452 16078 24454
rect 16210 32000 16266 32056
rect 15782 23418 15838 23420
rect 15862 23418 15918 23420
rect 15942 23418 15998 23420
rect 16022 23418 16078 23420
rect 15782 23366 15828 23418
rect 15828 23366 15838 23418
rect 15862 23366 15892 23418
rect 15892 23366 15904 23418
rect 15904 23366 15918 23418
rect 15942 23366 15956 23418
rect 15956 23366 15968 23418
rect 15968 23366 15998 23418
rect 16022 23366 16032 23418
rect 16032 23366 16078 23418
rect 15782 23364 15838 23366
rect 15862 23364 15918 23366
rect 15942 23364 15998 23366
rect 16022 23364 16078 23366
rect 15782 22330 15838 22332
rect 15862 22330 15918 22332
rect 15942 22330 15998 22332
rect 16022 22330 16078 22332
rect 15782 22278 15828 22330
rect 15828 22278 15838 22330
rect 15862 22278 15892 22330
rect 15892 22278 15904 22330
rect 15904 22278 15918 22330
rect 15942 22278 15956 22330
rect 15956 22278 15968 22330
rect 15968 22278 15998 22330
rect 16022 22278 16032 22330
rect 16032 22278 16078 22330
rect 15782 22276 15838 22278
rect 15862 22276 15918 22278
rect 15942 22276 15998 22278
rect 16022 22276 16078 22278
rect 15782 21242 15838 21244
rect 15862 21242 15918 21244
rect 15942 21242 15998 21244
rect 16022 21242 16078 21244
rect 15782 21190 15828 21242
rect 15828 21190 15838 21242
rect 15862 21190 15892 21242
rect 15892 21190 15904 21242
rect 15904 21190 15918 21242
rect 15942 21190 15956 21242
rect 15956 21190 15968 21242
rect 15968 21190 15998 21242
rect 16022 21190 16032 21242
rect 16032 21190 16078 21242
rect 15782 21188 15838 21190
rect 15862 21188 15918 21190
rect 15942 21188 15998 21190
rect 16022 21188 16078 21190
rect 16210 23160 16266 23216
rect 15782 20154 15838 20156
rect 15862 20154 15918 20156
rect 15942 20154 15998 20156
rect 16022 20154 16078 20156
rect 15782 20102 15828 20154
rect 15828 20102 15838 20154
rect 15862 20102 15892 20154
rect 15892 20102 15904 20154
rect 15904 20102 15918 20154
rect 15942 20102 15956 20154
rect 15956 20102 15968 20154
rect 15968 20102 15998 20154
rect 16022 20102 16032 20154
rect 16032 20102 16078 20154
rect 15782 20100 15838 20102
rect 15862 20100 15918 20102
rect 15942 20100 15998 20102
rect 16022 20100 16078 20102
rect 15782 19066 15838 19068
rect 15862 19066 15918 19068
rect 15942 19066 15998 19068
rect 16022 19066 16078 19068
rect 15782 19014 15828 19066
rect 15828 19014 15838 19066
rect 15862 19014 15892 19066
rect 15892 19014 15904 19066
rect 15904 19014 15918 19066
rect 15942 19014 15956 19066
rect 15956 19014 15968 19066
rect 15968 19014 15998 19066
rect 16022 19014 16032 19066
rect 16032 19014 16078 19066
rect 15782 19012 15838 19014
rect 15862 19012 15918 19014
rect 15942 19012 15998 19014
rect 16022 19012 16078 19014
rect 15782 17978 15838 17980
rect 15862 17978 15918 17980
rect 15942 17978 15998 17980
rect 16022 17978 16078 17980
rect 15782 17926 15828 17978
rect 15828 17926 15838 17978
rect 15862 17926 15892 17978
rect 15892 17926 15904 17978
rect 15904 17926 15918 17978
rect 15942 17926 15956 17978
rect 15956 17926 15968 17978
rect 15968 17926 15998 17978
rect 16022 17926 16032 17978
rect 16032 17926 16078 17978
rect 15782 17924 15838 17926
rect 15862 17924 15918 17926
rect 15942 17924 15998 17926
rect 16022 17924 16078 17926
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15942 16890 15998 16892
rect 16022 16890 16078 16892
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15904 16890
rect 15904 16838 15918 16890
rect 15942 16838 15956 16890
rect 15956 16838 15968 16890
rect 15968 16838 15998 16890
rect 16022 16838 16032 16890
rect 16032 16838 16078 16890
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 15942 16836 15998 16838
rect 16022 16836 16078 16838
rect 12817 11994 12873 11996
rect 12897 11994 12953 11996
rect 12977 11994 13033 11996
rect 13057 11994 13113 11996
rect 12817 11942 12863 11994
rect 12863 11942 12873 11994
rect 12897 11942 12927 11994
rect 12927 11942 12939 11994
rect 12939 11942 12953 11994
rect 12977 11942 12991 11994
rect 12991 11942 13003 11994
rect 13003 11942 13033 11994
rect 13057 11942 13067 11994
rect 13067 11942 13113 11994
rect 12817 11940 12873 11942
rect 12897 11940 12953 11942
rect 12977 11940 13033 11942
rect 13057 11940 13113 11942
rect 12817 10906 12873 10908
rect 12897 10906 12953 10908
rect 12977 10906 13033 10908
rect 13057 10906 13113 10908
rect 12817 10854 12863 10906
rect 12863 10854 12873 10906
rect 12897 10854 12927 10906
rect 12927 10854 12939 10906
rect 12939 10854 12953 10906
rect 12977 10854 12991 10906
rect 12991 10854 13003 10906
rect 13003 10854 13033 10906
rect 13057 10854 13067 10906
rect 13067 10854 13113 10906
rect 12817 10852 12873 10854
rect 12897 10852 12953 10854
rect 12977 10852 13033 10854
rect 13057 10852 13113 10854
rect 12817 9818 12873 9820
rect 12897 9818 12953 9820
rect 12977 9818 13033 9820
rect 13057 9818 13113 9820
rect 12817 9766 12863 9818
rect 12863 9766 12873 9818
rect 12897 9766 12927 9818
rect 12927 9766 12939 9818
rect 12939 9766 12953 9818
rect 12977 9766 12991 9818
rect 12991 9766 13003 9818
rect 13003 9766 13033 9818
rect 13057 9766 13067 9818
rect 13067 9766 13113 9818
rect 12817 9764 12873 9766
rect 12897 9764 12953 9766
rect 12977 9764 13033 9766
rect 13057 9764 13113 9766
rect 12817 8730 12873 8732
rect 12897 8730 12953 8732
rect 12977 8730 13033 8732
rect 13057 8730 13113 8732
rect 12817 8678 12863 8730
rect 12863 8678 12873 8730
rect 12897 8678 12927 8730
rect 12927 8678 12939 8730
rect 12939 8678 12953 8730
rect 12977 8678 12991 8730
rect 12991 8678 13003 8730
rect 13003 8678 13033 8730
rect 13057 8678 13067 8730
rect 13067 8678 13113 8730
rect 12817 8676 12873 8678
rect 12897 8676 12953 8678
rect 12977 8676 13033 8678
rect 13057 8676 13113 8678
rect 12817 7642 12873 7644
rect 12897 7642 12953 7644
rect 12977 7642 13033 7644
rect 13057 7642 13113 7644
rect 12817 7590 12863 7642
rect 12863 7590 12873 7642
rect 12897 7590 12927 7642
rect 12927 7590 12939 7642
rect 12939 7590 12953 7642
rect 12977 7590 12991 7642
rect 12991 7590 13003 7642
rect 13003 7590 13033 7642
rect 13057 7590 13067 7642
rect 13067 7590 13113 7642
rect 12817 7588 12873 7590
rect 12897 7588 12953 7590
rect 12977 7588 13033 7590
rect 13057 7588 13113 7590
rect 12817 6554 12873 6556
rect 12897 6554 12953 6556
rect 12977 6554 13033 6556
rect 13057 6554 13113 6556
rect 12817 6502 12863 6554
rect 12863 6502 12873 6554
rect 12897 6502 12927 6554
rect 12927 6502 12939 6554
rect 12939 6502 12953 6554
rect 12977 6502 12991 6554
rect 12991 6502 13003 6554
rect 13003 6502 13033 6554
rect 13057 6502 13067 6554
rect 13067 6502 13113 6554
rect 12817 6500 12873 6502
rect 12897 6500 12953 6502
rect 12977 6500 13033 6502
rect 13057 6500 13113 6502
rect 12817 5466 12873 5468
rect 12897 5466 12953 5468
rect 12977 5466 13033 5468
rect 13057 5466 13113 5468
rect 12817 5414 12863 5466
rect 12863 5414 12873 5466
rect 12897 5414 12927 5466
rect 12927 5414 12939 5466
rect 12939 5414 12953 5466
rect 12977 5414 12991 5466
rect 12991 5414 13003 5466
rect 13003 5414 13033 5466
rect 13057 5414 13067 5466
rect 13067 5414 13113 5466
rect 12817 5412 12873 5414
rect 12897 5412 12953 5414
rect 12977 5412 13033 5414
rect 13057 5412 13113 5414
rect 12817 4378 12873 4380
rect 12897 4378 12953 4380
rect 12977 4378 13033 4380
rect 13057 4378 13113 4380
rect 12817 4326 12863 4378
rect 12863 4326 12873 4378
rect 12897 4326 12927 4378
rect 12927 4326 12939 4378
rect 12939 4326 12953 4378
rect 12977 4326 12991 4378
rect 12991 4326 13003 4378
rect 13003 4326 13033 4378
rect 13057 4326 13067 4378
rect 13067 4326 13113 4378
rect 12817 4324 12873 4326
rect 12897 4324 12953 4326
rect 12977 4324 13033 4326
rect 13057 4324 13113 4326
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15942 15802 15998 15804
rect 16022 15802 16078 15804
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15904 15802
rect 15904 15750 15918 15802
rect 15942 15750 15956 15802
rect 15956 15750 15968 15802
rect 15968 15750 15998 15802
rect 16022 15750 16032 15802
rect 16032 15750 16078 15802
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 15942 15748 15998 15750
rect 16022 15748 16078 15750
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15942 14714 15998 14716
rect 16022 14714 16078 14716
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15904 14714
rect 15904 14662 15918 14714
rect 15942 14662 15956 14714
rect 15956 14662 15968 14714
rect 15968 14662 15998 14714
rect 16022 14662 16032 14714
rect 16032 14662 16078 14714
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 15942 14660 15998 14662
rect 16022 14660 16078 14662
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15942 13626 15998 13628
rect 16022 13626 16078 13628
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15904 13626
rect 15904 13574 15918 13626
rect 15942 13574 15956 13626
rect 15956 13574 15968 13626
rect 15968 13574 15998 13626
rect 16022 13574 16032 13626
rect 16032 13574 16078 13626
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15942 13572 15998 13574
rect 16022 13572 16078 13574
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15942 12538 15998 12540
rect 16022 12538 16078 12540
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15904 12538
rect 15904 12486 15918 12538
rect 15942 12486 15956 12538
rect 15956 12486 15968 12538
rect 15968 12486 15998 12538
rect 16022 12486 16032 12538
rect 16032 12486 16078 12538
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15942 12484 15998 12486
rect 16022 12484 16078 12486
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15942 11450 15998 11452
rect 16022 11450 16078 11452
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15904 11450
rect 15904 11398 15918 11450
rect 15942 11398 15956 11450
rect 15956 11398 15968 11450
rect 15968 11398 15998 11450
rect 16022 11398 16032 11450
rect 16032 11398 16078 11450
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 15942 11396 15998 11398
rect 16022 11396 16078 11398
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15942 10362 15998 10364
rect 16022 10362 16078 10364
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15904 10362
rect 15904 10310 15918 10362
rect 15942 10310 15956 10362
rect 15956 10310 15968 10362
rect 15968 10310 15998 10362
rect 16022 10310 16032 10362
rect 16032 10310 16078 10362
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 15942 10308 15998 10310
rect 16022 10308 16078 10310
rect 18142 14356 18144 14376
rect 18144 14356 18196 14376
rect 18196 14356 18198 14376
rect 18142 14320 18198 14356
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15942 9274 15998 9276
rect 16022 9274 16078 9276
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15904 9274
rect 15904 9222 15918 9274
rect 15942 9222 15956 9274
rect 15956 9222 15968 9274
rect 15968 9222 15998 9274
rect 16022 9222 16032 9274
rect 16032 9222 16078 9274
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 15942 9220 15998 9222
rect 16022 9220 16078 9222
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15942 8186 15998 8188
rect 16022 8186 16078 8188
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15904 8186
rect 15904 8134 15918 8186
rect 15942 8134 15956 8186
rect 15956 8134 15968 8186
rect 15968 8134 15998 8186
rect 16022 8134 16032 8186
rect 16032 8134 16078 8186
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15942 8132 15998 8134
rect 16022 8132 16078 8134
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15942 7098 15998 7100
rect 16022 7098 16078 7100
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15904 7098
rect 15904 7046 15918 7098
rect 15942 7046 15956 7098
rect 15956 7046 15968 7098
rect 15968 7046 15998 7098
rect 16022 7046 16032 7098
rect 16032 7046 16078 7098
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 15942 7044 15998 7046
rect 16022 7044 16078 7046
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15942 6010 15998 6012
rect 16022 6010 16078 6012
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15904 6010
rect 15904 5958 15918 6010
rect 15942 5958 15956 6010
rect 15956 5958 15968 6010
rect 15968 5958 15998 6010
rect 16022 5958 16032 6010
rect 16032 5958 16078 6010
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 15942 5956 15998 5958
rect 16022 5956 16078 5958
rect 17866 5480 17922 5536
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15942 4922 15998 4924
rect 16022 4922 16078 4924
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15904 4922
rect 15904 4870 15918 4922
rect 15942 4870 15956 4922
rect 15956 4870 15968 4922
rect 15968 4870 15998 4922
rect 16022 4870 16032 4922
rect 16032 4870 16078 4922
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 15942 4868 15998 4870
rect 16022 4868 16078 4870
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15942 3834 15998 3836
rect 16022 3834 16078 3836
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15904 3834
rect 15904 3782 15918 3834
rect 15942 3782 15956 3834
rect 15956 3782 15968 3834
rect 15968 3782 15998 3834
rect 16022 3782 16032 3834
rect 16032 3782 16078 3834
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 15942 3780 15998 3782
rect 16022 3780 16078 3782
rect 6886 3290 6942 3292
rect 6966 3290 7022 3292
rect 7046 3290 7102 3292
rect 7126 3290 7182 3292
rect 6886 3238 6932 3290
rect 6932 3238 6942 3290
rect 6966 3238 6996 3290
rect 6996 3238 7008 3290
rect 7008 3238 7022 3290
rect 7046 3238 7060 3290
rect 7060 3238 7072 3290
rect 7072 3238 7102 3290
rect 7126 3238 7136 3290
rect 7136 3238 7182 3290
rect 6886 3236 6942 3238
rect 6966 3236 7022 3238
rect 7046 3236 7102 3238
rect 7126 3236 7182 3238
rect 3921 2746 3977 2748
rect 4001 2746 4057 2748
rect 4081 2746 4137 2748
rect 4161 2746 4217 2748
rect 3921 2694 3967 2746
rect 3967 2694 3977 2746
rect 4001 2694 4031 2746
rect 4031 2694 4043 2746
rect 4043 2694 4057 2746
rect 4081 2694 4095 2746
rect 4095 2694 4107 2746
rect 4107 2694 4137 2746
rect 4161 2694 4171 2746
rect 4171 2694 4217 2746
rect 3921 2692 3977 2694
rect 4001 2692 4057 2694
rect 4081 2692 4137 2694
rect 4161 2692 4217 2694
rect 12817 3290 12873 3292
rect 12897 3290 12953 3292
rect 12977 3290 13033 3292
rect 13057 3290 13113 3292
rect 12817 3238 12863 3290
rect 12863 3238 12873 3290
rect 12897 3238 12927 3290
rect 12927 3238 12939 3290
rect 12939 3238 12953 3290
rect 12977 3238 12991 3290
rect 12991 3238 13003 3290
rect 13003 3238 13033 3290
rect 13057 3238 13067 3290
rect 13067 3238 13113 3290
rect 12817 3236 12873 3238
rect 12897 3236 12953 3238
rect 12977 3236 13033 3238
rect 13057 3236 13113 3238
rect 9852 2746 9908 2748
rect 9932 2746 9988 2748
rect 10012 2746 10068 2748
rect 10092 2746 10148 2748
rect 9852 2694 9898 2746
rect 9898 2694 9908 2746
rect 9932 2694 9962 2746
rect 9962 2694 9974 2746
rect 9974 2694 9988 2746
rect 10012 2694 10026 2746
rect 10026 2694 10038 2746
rect 10038 2694 10068 2746
rect 10092 2694 10102 2746
rect 10102 2694 10148 2746
rect 9852 2692 9908 2694
rect 9932 2692 9988 2694
rect 10012 2692 10068 2694
rect 10092 2692 10148 2694
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15942 2746 15998 2748
rect 16022 2746 16078 2748
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15904 2746
rect 15904 2694 15918 2746
rect 15942 2694 15956 2746
rect 15956 2694 15968 2746
rect 15968 2694 15998 2746
rect 16022 2694 16032 2746
rect 16032 2694 16078 2746
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 15942 2692 15998 2694
rect 16022 2692 16078 2694
rect 6886 2202 6942 2204
rect 6966 2202 7022 2204
rect 7046 2202 7102 2204
rect 7126 2202 7182 2204
rect 6886 2150 6932 2202
rect 6932 2150 6942 2202
rect 6966 2150 6996 2202
rect 6996 2150 7008 2202
rect 7008 2150 7022 2202
rect 7046 2150 7060 2202
rect 7060 2150 7072 2202
rect 7072 2150 7102 2202
rect 7126 2150 7136 2202
rect 7136 2150 7182 2202
rect 6886 2148 6942 2150
rect 6966 2148 7022 2150
rect 7046 2148 7102 2150
rect 7126 2148 7182 2150
rect 12817 2202 12873 2204
rect 12897 2202 12953 2204
rect 12977 2202 13033 2204
rect 13057 2202 13113 2204
rect 12817 2150 12863 2202
rect 12863 2150 12873 2202
rect 12897 2150 12927 2202
rect 12927 2150 12939 2202
rect 12939 2150 12953 2202
rect 12977 2150 12991 2202
rect 12991 2150 13003 2202
rect 13003 2150 13033 2202
rect 13057 2150 13067 2202
rect 13067 2150 13113 2202
rect 12817 2148 12873 2150
rect 12897 2148 12953 2150
rect 12977 2148 13033 2150
rect 13057 2148 13113 2150
<< metal3 >>
rect 3909 47360 4229 47361
rect 3909 47296 3917 47360
rect 3981 47296 3997 47360
rect 4061 47296 4077 47360
rect 4141 47296 4157 47360
rect 4221 47296 4229 47360
rect 3909 47295 4229 47296
rect 9840 47360 10160 47361
rect 9840 47296 9848 47360
rect 9912 47296 9928 47360
rect 9992 47296 10008 47360
rect 10072 47296 10088 47360
rect 10152 47296 10160 47360
rect 9840 47295 10160 47296
rect 15770 47360 16090 47361
rect 15770 47296 15778 47360
rect 15842 47296 15858 47360
rect 15922 47296 15938 47360
rect 16002 47296 16018 47360
rect 16082 47296 16090 47360
rect 15770 47295 16090 47296
rect 6874 46816 7194 46817
rect 6874 46752 6882 46816
rect 6946 46752 6962 46816
rect 7026 46752 7042 46816
rect 7106 46752 7122 46816
rect 7186 46752 7194 46816
rect 6874 46751 7194 46752
rect 12805 46816 13125 46817
rect 12805 46752 12813 46816
rect 12877 46752 12893 46816
rect 12957 46752 12973 46816
rect 13037 46752 13053 46816
rect 13117 46752 13125 46816
rect 12805 46751 13125 46752
rect 3909 46272 4229 46273
rect 3909 46208 3917 46272
rect 3981 46208 3997 46272
rect 4061 46208 4077 46272
rect 4141 46208 4157 46272
rect 4221 46208 4229 46272
rect 3909 46207 4229 46208
rect 9840 46272 10160 46273
rect 9840 46208 9848 46272
rect 9912 46208 9928 46272
rect 9992 46208 10008 46272
rect 10072 46208 10088 46272
rect 10152 46208 10160 46272
rect 9840 46207 10160 46208
rect 15770 46272 16090 46273
rect 15770 46208 15778 46272
rect 15842 46208 15858 46272
rect 15922 46208 15938 46272
rect 16002 46208 16018 46272
rect 16082 46208 16090 46272
rect 15770 46207 16090 46208
rect 6874 45728 7194 45729
rect 6874 45664 6882 45728
rect 6946 45664 6962 45728
rect 7026 45664 7042 45728
rect 7106 45664 7122 45728
rect 7186 45664 7194 45728
rect 6874 45663 7194 45664
rect 12805 45728 13125 45729
rect 12805 45664 12813 45728
rect 12877 45664 12893 45728
rect 12957 45664 12973 45728
rect 13037 45664 13053 45728
rect 13117 45664 13125 45728
rect 12805 45663 13125 45664
rect 3909 45184 4229 45185
rect 3909 45120 3917 45184
rect 3981 45120 3997 45184
rect 4061 45120 4077 45184
rect 4141 45120 4157 45184
rect 4221 45120 4229 45184
rect 3909 45119 4229 45120
rect 9840 45184 10160 45185
rect 9840 45120 9848 45184
rect 9912 45120 9928 45184
rect 9992 45120 10008 45184
rect 10072 45120 10088 45184
rect 10152 45120 10160 45184
rect 9840 45119 10160 45120
rect 15770 45184 16090 45185
rect 15770 45120 15778 45184
rect 15842 45120 15858 45184
rect 15922 45120 15938 45184
rect 16002 45120 16018 45184
rect 16082 45120 16090 45184
rect 15770 45119 16090 45120
rect 6874 44640 7194 44641
rect 6874 44576 6882 44640
rect 6946 44576 6962 44640
rect 7026 44576 7042 44640
rect 7106 44576 7122 44640
rect 7186 44576 7194 44640
rect 6874 44575 7194 44576
rect 12805 44640 13125 44641
rect 12805 44576 12813 44640
rect 12877 44576 12893 44640
rect 12957 44576 12973 44640
rect 13037 44576 13053 44640
rect 13117 44576 13125 44640
rect 12805 44575 13125 44576
rect 0 44298 800 44328
rect 1853 44298 1919 44301
rect 0 44296 1919 44298
rect 0 44240 1858 44296
rect 1914 44240 1919 44296
rect 0 44238 1919 44240
rect 0 44208 800 44238
rect 1853 44235 1919 44238
rect 3909 44096 4229 44097
rect 3909 44032 3917 44096
rect 3981 44032 3997 44096
rect 4061 44032 4077 44096
rect 4141 44032 4157 44096
rect 4221 44032 4229 44096
rect 3909 44031 4229 44032
rect 9840 44096 10160 44097
rect 9840 44032 9848 44096
rect 9912 44032 9928 44096
rect 9992 44032 10008 44096
rect 10072 44032 10088 44096
rect 10152 44032 10160 44096
rect 9840 44031 10160 44032
rect 15770 44096 16090 44097
rect 15770 44032 15778 44096
rect 15842 44032 15858 44096
rect 15922 44032 15938 44096
rect 16002 44032 16018 44096
rect 16082 44032 16090 44096
rect 15770 44031 16090 44032
rect 6874 43552 7194 43553
rect 6874 43488 6882 43552
rect 6946 43488 6962 43552
rect 7026 43488 7042 43552
rect 7106 43488 7122 43552
rect 7186 43488 7194 43552
rect 6874 43487 7194 43488
rect 12805 43552 13125 43553
rect 12805 43488 12813 43552
rect 12877 43488 12893 43552
rect 12957 43488 12973 43552
rect 13037 43488 13053 43552
rect 13117 43488 13125 43552
rect 12805 43487 13125 43488
rect 3909 43008 4229 43009
rect 3909 42944 3917 43008
rect 3981 42944 3997 43008
rect 4061 42944 4077 43008
rect 4141 42944 4157 43008
rect 4221 42944 4229 43008
rect 3909 42943 4229 42944
rect 9840 43008 10160 43009
rect 9840 42944 9848 43008
rect 9912 42944 9928 43008
rect 9992 42944 10008 43008
rect 10072 42944 10088 43008
rect 10152 42944 10160 43008
rect 9840 42943 10160 42944
rect 15770 43008 16090 43009
rect 15770 42944 15778 43008
rect 15842 42944 15858 43008
rect 15922 42944 15938 43008
rect 16002 42944 16018 43008
rect 16082 42944 16090 43008
rect 15770 42943 16090 42944
rect 6874 42464 7194 42465
rect 6874 42400 6882 42464
rect 6946 42400 6962 42464
rect 7026 42400 7042 42464
rect 7106 42400 7122 42464
rect 7186 42400 7194 42464
rect 6874 42399 7194 42400
rect 12805 42464 13125 42465
rect 12805 42400 12813 42464
rect 12877 42400 12893 42464
rect 12957 42400 12973 42464
rect 13037 42400 13053 42464
rect 13117 42400 13125 42464
rect 12805 42399 13125 42400
rect 3909 41920 4229 41921
rect 3909 41856 3917 41920
rect 3981 41856 3997 41920
rect 4061 41856 4077 41920
rect 4141 41856 4157 41920
rect 4221 41856 4229 41920
rect 3909 41855 4229 41856
rect 9840 41920 10160 41921
rect 9840 41856 9848 41920
rect 9912 41856 9928 41920
rect 9992 41856 10008 41920
rect 10072 41856 10088 41920
rect 10152 41856 10160 41920
rect 9840 41855 10160 41856
rect 15770 41920 16090 41921
rect 15770 41856 15778 41920
rect 15842 41856 15858 41920
rect 15922 41856 15938 41920
rect 16002 41856 16018 41920
rect 16082 41856 16090 41920
rect 15770 41855 16090 41856
rect 6874 41376 7194 41377
rect 6874 41312 6882 41376
rect 6946 41312 6962 41376
rect 7026 41312 7042 41376
rect 7106 41312 7122 41376
rect 7186 41312 7194 41376
rect 6874 41311 7194 41312
rect 12805 41376 13125 41377
rect 12805 41312 12813 41376
rect 12877 41312 12893 41376
rect 12957 41312 12973 41376
rect 13037 41312 13053 41376
rect 13117 41312 13125 41376
rect 12805 41311 13125 41312
rect 18137 40898 18203 40901
rect 19200 40898 20000 40928
rect 18137 40896 20000 40898
rect 18137 40840 18142 40896
rect 18198 40840 20000 40896
rect 18137 40838 20000 40840
rect 18137 40835 18203 40838
rect 3909 40832 4229 40833
rect 3909 40768 3917 40832
rect 3981 40768 3997 40832
rect 4061 40768 4077 40832
rect 4141 40768 4157 40832
rect 4221 40768 4229 40832
rect 3909 40767 4229 40768
rect 9840 40832 10160 40833
rect 9840 40768 9848 40832
rect 9912 40768 9928 40832
rect 9992 40768 10008 40832
rect 10072 40768 10088 40832
rect 10152 40768 10160 40832
rect 9840 40767 10160 40768
rect 15770 40832 16090 40833
rect 15770 40768 15778 40832
rect 15842 40768 15858 40832
rect 15922 40768 15938 40832
rect 16002 40768 16018 40832
rect 16082 40768 16090 40832
rect 19200 40808 20000 40838
rect 15770 40767 16090 40768
rect 6874 40288 7194 40289
rect 6874 40224 6882 40288
rect 6946 40224 6962 40288
rect 7026 40224 7042 40288
rect 7106 40224 7122 40288
rect 7186 40224 7194 40288
rect 6874 40223 7194 40224
rect 12805 40288 13125 40289
rect 12805 40224 12813 40288
rect 12877 40224 12893 40288
rect 12957 40224 12973 40288
rect 13037 40224 13053 40288
rect 13117 40224 13125 40288
rect 12805 40223 13125 40224
rect 3909 39744 4229 39745
rect 3909 39680 3917 39744
rect 3981 39680 3997 39744
rect 4061 39680 4077 39744
rect 4141 39680 4157 39744
rect 4221 39680 4229 39744
rect 3909 39679 4229 39680
rect 9840 39744 10160 39745
rect 9840 39680 9848 39744
rect 9912 39680 9928 39744
rect 9992 39680 10008 39744
rect 10072 39680 10088 39744
rect 10152 39680 10160 39744
rect 9840 39679 10160 39680
rect 15770 39744 16090 39745
rect 15770 39680 15778 39744
rect 15842 39680 15858 39744
rect 15922 39680 15938 39744
rect 16002 39680 16018 39744
rect 16082 39680 16090 39744
rect 15770 39679 16090 39680
rect 6874 39200 7194 39201
rect 6874 39136 6882 39200
rect 6946 39136 6962 39200
rect 7026 39136 7042 39200
rect 7106 39136 7122 39200
rect 7186 39136 7194 39200
rect 6874 39135 7194 39136
rect 12805 39200 13125 39201
rect 12805 39136 12813 39200
rect 12877 39136 12893 39200
rect 12957 39136 12973 39200
rect 13037 39136 13053 39200
rect 13117 39136 13125 39200
rect 12805 39135 13125 39136
rect 3909 38656 4229 38657
rect 3909 38592 3917 38656
rect 3981 38592 3997 38656
rect 4061 38592 4077 38656
rect 4141 38592 4157 38656
rect 4221 38592 4229 38656
rect 3909 38591 4229 38592
rect 9840 38656 10160 38657
rect 9840 38592 9848 38656
rect 9912 38592 9928 38656
rect 9992 38592 10008 38656
rect 10072 38592 10088 38656
rect 10152 38592 10160 38656
rect 9840 38591 10160 38592
rect 15770 38656 16090 38657
rect 15770 38592 15778 38656
rect 15842 38592 15858 38656
rect 15922 38592 15938 38656
rect 16002 38592 16018 38656
rect 16082 38592 16090 38656
rect 15770 38591 16090 38592
rect 6874 38112 7194 38113
rect 6874 38048 6882 38112
rect 6946 38048 6962 38112
rect 7026 38048 7042 38112
rect 7106 38048 7122 38112
rect 7186 38048 7194 38112
rect 6874 38047 7194 38048
rect 12805 38112 13125 38113
rect 12805 38048 12813 38112
rect 12877 38048 12893 38112
rect 12957 38048 12973 38112
rect 13037 38048 13053 38112
rect 13117 38048 13125 38112
rect 12805 38047 13125 38048
rect 3909 37568 4229 37569
rect 3909 37504 3917 37568
rect 3981 37504 3997 37568
rect 4061 37504 4077 37568
rect 4141 37504 4157 37568
rect 4221 37504 4229 37568
rect 3909 37503 4229 37504
rect 9840 37568 10160 37569
rect 9840 37504 9848 37568
rect 9912 37504 9928 37568
rect 9992 37504 10008 37568
rect 10072 37504 10088 37568
rect 10152 37504 10160 37568
rect 9840 37503 10160 37504
rect 15770 37568 16090 37569
rect 15770 37504 15778 37568
rect 15842 37504 15858 37568
rect 15922 37504 15938 37568
rect 16002 37504 16018 37568
rect 16082 37504 16090 37568
rect 15770 37503 16090 37504
rect 6874 37024 7194 37025
rect 6874 36960 6882 37024
rect 6946 36960 6962 37024
rect 7026 36960 7042 37024
rect 7106 36960 7122 37024
rect 7186 36960 7194 37024
rect 6874 36959 7194 36960
rect 12805 37024 13125 37025
rect 12805 36960 12813 37024
rect 12877 36960 12893 37024
rect 12957 36960 12973 37024
rect 13037 36960 13053 37024
rect 13117 36960 13125 37024
rect 12805 36959 13125 36960
rect 3909 36480 4229 36481
rect 3909 36416 3917 36480
rect 3981 36416 3997 36480
rect 4061 36416 4077 36480
rect 4141 36416 4157 36480
rect 4221 36416 4229 36480
rect 3909 36415 4229 36416
rect 9840 36480 10160 36481
rect 9840 36416 9848 36480
rect 9912 36416 9928 36480
rect 9992 36416 10008 36480
rect 10072 36416 10088 36480
rect 10152 36416 10160 36480
rect 9840 36415 10160 36416
rect 15770 36480 16090 36481
rect 15770 36416 15778 36480
rect 15842 36416 15858 36480
rect 15922 36416 15938 36480
rect 16002 36416 16018 36480
rect 16082 36416 16090 36480
rect 15770 36415 16090 36416
rect 6874 35936 7194 35937
rect 6874 35872 6882 35936
rect 6946 35872 6962 35936
rect 7026 35872 7042 35936
rect 7106 35872 7122 35936
rect 7186 35872 7194 35936
rect 6874 35871 7194 35872
rect 12805 35936 13125 35937
rect 12805 35872 12813 35936
rect 12877 35872 12893 35936
rect 12957 35872 12973 35936
rect 13037 35872 13053 35936
rect 13117 35872 13125 35936
rect 12805 35871 13125 35872
rect 0 35458 800 35488
rect 1393 35458 1459 35461
rect 0 35456 1459 35458
rect 0 35400 1398 35456
rect 1454 35400 1459 35456
rect 0 35398 1459 35400
rect 0 35368 800 35398
rect 1393 35395 1459 35398
rect 3909 35392 4229 35393
rect 3909 35328 3917 35392
rect 3981 35328 3997 35392
rect 4061 35328 4077 35392
rect 4141 35328 4157 35392
rect 4221 35328 4229 35392
rect 3909 35327 4229 35328
rect 9840 35392 10160 35393
rect 9840 35328 9848 35392
rect 9912 35328 9928 35392
rect 9992 35328 10008 35392
rect 10072 35328 10088 35392
rect 10152 35328 10160 35392
rect 9840 35327 10160 35328
rect 15770 35392 16090 35393
rect 15770 35328 15778 35392
rect 15842 35328 15858 35392
rect 15922 35328 15938 35392
rect 16002 35328 16018 35392
rect 16082 35328 16090 35392
rect 15770 35327 16090 35328
rect 6874 34848 7194 34849
rect 6874 34784 6882 34848
rect 6946 34784 6962 34848
rect 7026 34784 7042 34848
rect 7106 34784 7122 34848
rect 7186 34784 7194 34848
rect 6874 34783 7194 34784
rect 12805 34848 13125 34849
rect 12805 34784 12813 34848
rect 12877 34784 12893 34848
rect 12957 34784 12973 34848
rect 13037 34784 13053 34848
rect 13117 34784 13125 34848
rect 12805 34783 13125 34784
rect 3909 34304 4229 34305
rect 3909 34240 3917 34304
rect 3981 34240 3997 34304
rect 4061 34240 4077 34304
rect 4141 34240 4157 34304
rect 4221 34240 4229 34304
rect 3909 34239 4229 34240
rect 9840 34304 10160 34305
rect 9840 34240 9848 34304
rect 9912 34240 9928 34304
rect 9992 34240 10008 34304
rect 10072 34240 10088 34304
rect 10152 34240 10160 34304
rect 9840 34239 10160 34240
rect 15770 34304 16090 34305
rect 15770 34240 15778 34304
rect 15842 34240 15858 34304
rect 15922 34240 15938 34304
rect 16002 34240 16018 34304
rect 16082 34240 16090 34304
rect 15770 34239 16090 34240
rect 6874 33760 7194 33761
rect 6874 33696 6882 33760
rect 6946 33696 6962 33760
rect 7026 33696 7042 33760
rect 7106 33696 7122 33760
rect 7186 33696 7194 33760
rect 6874 33695 7194 33696
rect 12805 33760 13125 33761
rect 12805 33696 12813 33760
rect 12877 33696 12893 33760
rect 12957 33696 12973 33760
rect 13037 33696 13053 33760
rect 13117 33696 13125 33760
rect 12805 33695 13125 33696
rect 3909 33216 4229 33217
rect 3909 33152 3917 33216
rect 3981 33152 3997 33216
rect 4061 33152 4077 33216
rect 4141 33152 4157 33216
rect 4221 33152 4229 33216
rect 3909 33151 4229 33152
rect 9840 33216 10160 33217
rect 9840 33152 9848 33216
rect 9912 33152 9928 33216
rect 9992 33152 10008 33216
rect 10072 33152 10088 33216
rect 10152 33152 10160 33216
rect 9840 33151 10160 33152
rect 15770 33216 16090 33217
rect 15770 33152 15778 33216
rect 15842 33152 15858 33216
rect 15922 33152 15938 33216
rect 16002 33152 16018 33216
rect 16082 33152 16090 33216
rect 15770 33151 16090 33152
rect 5993 33146 6059 33149
rect 7925 33146 7991 33149
rect 5993 33144 7991 33146
rect 5993 33088 5998 33144
rect 6054 33088 7930 33144
rect 7986 33088 7991 33144
rect 5993 33086 7991 33088
rect 5993 33083 6059 33086
rect 7925 33083 7991 33086
rect 6874 32672 7194 32673
rect 6874 32608 6882 32672
rect 6946 32608 6962 32672
rect 7026 32608 7042 32672
rect 7106 32608 7122 32672
rect 7186 32608 7194 32672
rect 6874 32607 7194 32608
rect 12805 32672 13125 32673
rect 12805 32608 12813 32672
rect 12877 32608 12893 32672
rect 12957 32608 12973 32672
rect 13037 32608 13053 32672
rect 13117 32608 13125 32672
rect 12805 32607 13125 32608
rect 3909 32128 4229 32129
rect 3909 32064 3917 32128
rect 3981 32064 3997 32128
rect 4061 32064 4077 32128
rect 4141 32064 4157 32128
rect 4221 32064 4229 32128
rect 3909 32063 4229 32064
rect 9840 32128 10160 32129
rect 9840 32064 9848 32128
rect 9912 32064 9928 32128
rect 9992 32064 10008 32128
rect 10072 32064 10088 32128
rect 10152 32064 10160 32128
rect 9840 32063 10160 32064
rect 15770 32128 16090 32129
rect 15770 32064 15778 32128
rect 15842 32064 15858 32128
rect 15922 32064 15938 32128
rect 16002 32064 16018 32128
rect 16082 32064 16090 32128
rect 15770 32063 16090 32064
rect 16205 32058 16271 32061
rect 19200 32058 20000 32088
rect 16205 32056 20000 32058
rect 16205 32000 16210 32056
rect 16266 32000 20000 32056
rect 16205 31998 20000 32000
rect 16205 31995 16271 31998
rect 19200 31968 20000 31998
rect 6874 31584 7194 31585
rect 6874 31520 6882 31584
rect 6946 31520 6962 31584
rect 7026 31520 7042 31584
rect 7106 31520 7122 31584
rect 7186 31520 7194 31584
rect 6874 31519 7194 31520
rect 12805 31584 13125 31585
rect 12805 31520 12813 31584
rect 12877 31520 12893 31584
rect 12957 31520 12973 31584
rect 13037 31520 13053 31584
rect 13117 31520 13125 31584
rect 12805 31519 13125 31520
rect 3909 31040 4229 31041
rect 3909 30976 3917 31040
rect 3981 30976 3997 31040
rect 4061 30976 4077 31040
rect 4141 30976 4157 31040
rect 4221 30976 4229 31040
rect 3909 30975 4229 30976
rect 9840 31040 10160 31041
rect 9840 30976 9848 31040
rect 9912 30976 9928 31040
rect 9992 30976 10008 31040
rect 10072 30976 10088 31040
rect 10152 30976 10160 31040
rect 9840 30975 10160 30976
rect 15770 31040 16090 31041
rect 15770 30976 15778 31040
rect 15842 30976 15858 31040
rect 15922 30976 15938 31040
rect 16002 30976 16018 31040
rect 16082 30976 16090 31040
rect 15770 30975 16090 30976
rect 6874 30496 7194 30497
rect 6874 30432 6882 30496
rect 6946 30432 6962 30496
rect 7026 30432 7042 30496
rect 7106 30432 7122 30496
rect 7186 30432 7194 30496
rect 6874 30431 7194 30432
rect 12805 30496 13125 30497
rect 12805 30432 12813 30496
rect 12877 30432 12893 30496
rect 12957 30432 12973 30496
rect 13037 30432 13053 30496
rect 13117 30432 13125 30496
rect 12805 30431 13125 30432
rect 3909 29952 4229 29953
rect 3909 29888 3917 29952
rect 3981 29888 3997 29952
rect 4061 29888 4077 29952
rect 4141 29888 4157 29952
rect 4221 29888 4229 29952
rect 3909 29887 4229 29888
rect 9840 29952 10160 29953
rect 9840 29888 9848 29952
rect 9912 29888 9928 29952
rect 9992 29888 10008 29952
rect 10072 29888 10088 29952
rect 10152 29888 10160 29952
rect 9840 29887 10160 29888
rect 15770 29952 16090 29953
rect 15770 29888 15778 29952
rect 15842 29888 15858 29952
rect 15922 29888 15938 29952
rect 16002 29888 16018 29952
rect 16082 29888 16090 29952
rect 15770 29887 16090 29888
rect 6874 29408 7194 29409
rect 6874 29344 6882 29408
rect 6946 29344 6962 29408
rect 7026 29344 7042 29408
rect 7106 29344 7122 29408
rect 7186 29344 7194 29408
rect 6874 29343 7194 29344
rect 12805 29408 13125 29409
rect 12805 29344 12813 29408
rect 12877 29344 12893 29408
rect 12957 29344 12973 29408
rect 13037 29344 13053 29408
rect 13117 29344 13125 29408
rect 12805 29343 13125 29344
rect 3909 28864 4229 28865
rect 3909 28800 3917 28864
rect 3981 28800 3997 28864
rect 4061 28800 4077 28864
rect 4141 28800 4157 28864
rect 4221 28800 4229 28864
rect 3909 28799 4229 28800
rect 9840 28864 10160 28865
rect 9840 28800 9848 28864
rect 9912 28800 9928 28864
rect 9992 28800 10008 28864
rect 10072 28800 10088 28864
rect 10152 28800 10160 28864
rect 9840 28799 10160 28800
rect 15770 28864 16090 28865
rect 15770 28800 15778 28864
rect 15842 28800 15858 28864
rect 15922 28800 15938 28864
rect 16002 28800 16018 28864
rect 16082 28800 16090 28864
rect 15770 28799 16090 28800
rect 6874 28320 7194 28321
rect 6874 28256 6882 28320
rect 6946 28256 6962 28320
rect 7026 28256 7042 28320
rect 7106 28256 7122 28320
rect 7186 28256 7194 28320
rect 6874 28255 7194 28256
rect 12805 28320 13125 28321
rect 12805 28256 12813 28320
rect 12877 28256 12893 28320
rect 12957 28256 12973 28320
rect 13037 28256 13053 28320
rect 13117 28256 13125 28320
rect 12805 28255 13125 28256
rect 3909 27776 4229 27777
rect 3909 27712 3917 27776
rect 3981 27712 3997 27776
rect 4061 27712 4077 27776
rect 4141 27712 4157 27776
rect 4221 27712 4229 27776
rect 3909 27711 4229 27712
rect 9840 27776 10160 27777
rect 9840 27712 9848 27776
rect 9912 27712 9928 27776
rect 9992 27712 10008 27776
rect 10072 27712 10088 27776
rect 10152 27712 10160 27776
rect 9840 27711 10160 27712
rect 15770 27776 16090 27777
rect 15770 27712 15778 27776
rect 15842 27712 15858 27776
rect 15922 27712 15938 27776
rect 16002 27712 16018 27776
rect 16082 27712 16090 27776
rect 15770 27711 16090 27712
rect 6874 27232 7194 27233
rect 6874 27168 6882 27232
rect 6946 27168 6962 27232
rect 7026 27168 7042 27232
rect 7106 27168 7122 27232
rect 7186 27168 7194 27232
rect 6874 27167 7194 27168
rect 12805 27232 13125 27233
rect 12805 27168 12813 27232
rect 12877 27168 12893 27232
rect 12957 27168 12973 27232
rect 13037 27168 13053 27232
rect 13117 27168 13125 27232
rect 12805 27167 13125 27168
rect 3909 26688 4229 26689
rect 0 26618 800 26648
rect 3909 26624 3917 26688
rect 3981 26624 3997 26688
rect 4061 26624 4077 26688
rect 4141 26624 4157 26688
rect 4221 26624 4229 26688
rect 3909 26623 4229 26624
rect 9840 26688 10160 26689
rect 9840 26624 9848 26688
rect 9912 26624 9928 26688
rect 9992 26624 10008 26688
rect 10072 26624 10088 26688
rect 10152 26624 10160 26688
rect 9840 26623 10160 26624
rect 15770 26688 16090 26689
rect 15770 26624 15778 26688
rect 15842 26624 15858 26688
rect 15922 26624 15938 26688
rect 16002 26624 16018 26688
rect 16082 26624 16090 26688
rect 15770 26623 16090 26624
rect 1485 26618 1551 26621
rect 0 26616 1551 26618
rect 0 26560 1490 26616
rect 1546 26560 1551 26616
rect 0 26558 1551 26560
rect 0 26528 800 26558
rect 1485 26555 1551 26558
rect 6874 26144 7194 26145
rect 6874 26080 6882 26144
rect 6946 26080 6962 26144
rect 7026 26080 7042 26144
rect 7106 26080 7122 26144
rect 7186 26080 7194 26144
rect 6874 26079 7194 26080
rect 12805 26144 13125 26145
rect 12805 26080 12813 26144
rect 12877 26080 12893 26144
rect 12957 26080 12973 26144
rect 13037 26080 13053 26144
rect 13117 26080 13125 26144
rect 12805 26079 13125 26080
rect 3909 25600 4229 25601
rect 3909 25536 3917 25600
rect 3981 25536 3997 25600
rect 4061 25536 4077 25600
rect 4141 25536 4157 25600
rect 4221 25536 4229 25600
rect 3909 25535 4229 25536
rect 9840 25600 10160 25601
rect 9840 25536 9848 25600
rect 9912 25536 9928 25600
rect 9992 25536 10008 25600
rect 10072 25536 10088 25600
rect 10152 25536 10160 25600
rect 9840 25535 10160 25536
rect 15770 25600 16090 25601
rect 15770 25536 15778 25600
rect 15842 25536 15858 25600
rect 15922 25536 15938 25600
rect 16002 25536 16018 25600
rect 16082 25536 16090 25600
rect 15770 25535 16090 25536
rect 6874 25056 7194 25057
rect 6874 24992 6882 25056
rect 6946 24992 6962 25056
rect 7026 24992 7042 25056
rect 7106 24992 7122 25056
rect 7186 24992 7194 25056
rect 6874 24991 7194 24992
rect 12805 25056 13125 25057
rect 12805 24992 12813 25056
rect 12877 24992 12893 25056
rect 12957 24992 12973 25056
rect 13037 24992 13053 25056
rect 13117 24992 13125 25056
rect 12805 24991 13125 24992
rect 3909 24512 4229 24513
rect 3909 24448 3917 24512
rect 3981 24448 3997 24512
rect 4061 24448 4077 24512
rect 4141 24448 4157 24512
rect 4221 24448 4229 24512
rect 3909 24447 4229 24448
rect 9840 24512 10160 24513
rect 9840 24448 9848 24512
rect 9912 24448 9928 24512
rect 9992 24448 10008 24512
rect 10072 24448 10088 24512
rect 10152 24448 10160 24512
rect 9840 24447 10160 24448
rect 15770 24512 16090 24513
rect 15770 24448 15778 24512
rect 15842 24448 15858 24512
rect 15922 24448 15938 24512
rect 16002 24448 16018 24512
rect 16082 24448 16090 24512
rect 15770 24447 16090 24448
rect 6874 23968 7194 23969
rect 6874 23904 6882 23968
rect 6946 23904 6962 23968
rect 7026 23904 7042 23968
rect 7106 23904 7122 23968
rect 7186 23904 7194 23968
rect 6874 23903 7194 23904
rect 12805 23968 13125 23969
rect 12805 23904 12813 23968
rect 12877 23904 12893 23968
rect 12957 23904 12973 23968
rect 13037 23904 13053 23968
rect 13117 23904 13125 23968
rect 12805 23903 13125 23904
rect 3909 23424 4229 23425
rect 3909 23360 3917 23424
rect 3981 23360 3997 23424
rect 4061 23360 4077 23424
rect 4141 23360 4157 23424
rect 4221 23360 4229 23424
rect 3909 23359 4229 23360
rect 9840 23424 10160 23425
rect 9840 23360 9848 23424
rect 9912 23360 9928 23424
rect 9992 23360 10008 23424
rect 10072 23360 10088 23424
rect 10152 23360 10160 23424
rect 9840 23359 10160 23360
rect 15770 23424 16090 23425
rect 15770 23360 15778 23424
rect 15842 23360 15858 23424
rect 15922 23360 15938 23424
rect 16002 23360 16018 23424
rect 16082 23360 16090 23424
rect 15770 23359 16090 23360
rect 16205 23218 16271 23221
rect 19200 23218 20000 23248
rect 16205 23216 20000 23218
rect 16205 23160 16210 23216
rect 16266 23160 20000 23216
rect 16205 23158 20000 23160
rect 16205 23155 16271 23158
rect 19200 23128 20000 23158
rect 6874 22880 7194 22881
rect 6874 22816 6882 22880
rect 6946 22816 6962 22880
rect 7026 22816 7042 22880
rect 7106 22816 7122 22880
rect 7186 22816 7194 22880
rect 6874 22815 7194 22816
rect 12805 22880 13125 22881
rect 12805 22816 12813 22880
rect 12877 22816 12893 22880
rect 12957 22816 12973 22880
rect 13037 22816 13053 22880
rect 13117 22816 13125 22880
rect 12805 22815 13125 22816
rect 3909 22336 4229 22337
rect 3909 22272 3917 22336
rect 3981 22272 3997 22336
rect 4061 22272 4077 22336
rect 4141 22272 4157 22336
rect 4221 22272 4229 22336
rect 3909 22271 4229 22272
rect 9840 22336 10160 22337
rect 9840 22272 9848 22336
rect 9912 22272 9928 22336
rect 9992 22272 10008 22336
rect 10072 22272 10088 22336
rect 10152 22272 10160 22336
rect 9840 22271 10160 22272
rect 15770 22336 16090 22337
rect 15770 22272 15778 22336
rect 15842 22272 15858 22336
rect 15922 22272 15938 22336
rect 16002 22272 16018 22336
rect 16082 22272 16090 22336
rect 15770 22271 16090 22272
rect 6874 21792 7194 21793
rect 6874 21728 6882 21792
rect 6946 21728 6962 21792
rect 7026 21728 7042 21792
rect 7106 21728 7122 21792
rect 7186 21728 7194 21792
rect 6874 21727 7194 21728
rect 12805 21792 13125 21793
rect 12805 21728 12813 21792
rect 12877 21728 12893 21792
rect 12957 21728 12973 21792
rect 13037 21728 13053 21792
rect 13117 21728 13125 21792
rect 12805 21727 13125 21728
rect 3909 21248 4229 21249
rect 3909 21184 3917 21248
rect 3981 21184 3997 21248
rect 4061 21184 4077 21248
rect 4141 21184 4157 21248
rect 4221 21184 4229 21248
rect 3909 21183 4229 21184
rect 9840 21248 10160 21249
rect 9840 21184 9848 21248
rect 9912 21184 9928 21248
rect 9992 21184 10008 21248
rect 10072 21184 10088 21248
rect 10152 21184 10160 21248
rect 9840 21183 10160 21184
rect 15770 21248 16090 21249
rect 15770 21184 15778 21248
rect 15842 21184 15858 21248
rect 15922 21184 15938 21248
rect 16002 21184 16018 21248
rect 16082 21184 16090 21248
rect 15770 21183 16090 21184
rect 6874 20704 7194 20705
rect 6874 20640 6882 20704
rect 6946 20640 6962 20704
rect 7026 20640 7042 20704
rect 7106 20640 7122 20704
rect 7186 20640 7194 20704
rect 6874 20639 7194 20640
rect 12805 20704 13125 20705
rect 12805 20640 12813 20704
rect 12877 20640 12893 20704
rect 12957 20640 12973 20704
rect 13037 20640 13053 20704
rect 13117 20640 13125 20704
rect 12805 20639 13125 20640
rect 3909 20160 4229 20161
rect 3909 20096 3917 20160
rect 3981 20096 3997 20160
rect 4061 20096 4077 20160
rect 4141 20096 4157 20160
rect 4221 20096 4229 20160
rect 3909 20095 4229 20096
rect 9840 20160 10160 20161
rect 9840 20096 9848 20160
rect 9912 20096 9928 20160
rect 9992 20096 10008 20160
rect 10072 20096 10088 20160
rect 10152 20096 10160 20160
rect 9840 20095 10160 20096
rect 15770 20160 16090 20161
rect 15770 20096 15778 20160
rect 15842 20096 15858 20160
rect 15922 20096 15938 20160
rect 16002 20096 16018 20160
rect 16082 20096 16090 20160
rect 15770 20095 16090 20096
rect 6874 19616 7194 19617
rect 6874 19552 6882 19616
rect 6946 19552 6962 19616
rect 7026 19552 7042 19616
rect 7106 19552 7122 19616
rect 7186 19552 7194 19616
rect 6874 19551 7194 19552
rect 12805 19616 13125 19617
rect 12805 19552 12813 19616
rect 12877 19552 12893 19616
rect 12957 19552 12973 19616
rect 13037 19552 13053 19616
rect 13117 19552 13125 19616
rect 12805 19551 13125 19552
rect 3909 19072 4229 19073
rect 3909 19008 3917 19072
rect 3981 19008 3997 19072
rect 4061 19008 4077 19072
rect 4141 19008 4157 19072
rect 4221 19008 4229 19072
rect 3909 19007 4229 19008
rect 9840 19072 10160 19073
rect 9840 19008 9848 19072
rect 9912 19008 9928 19072
rect 9992 19008 10008 19072
rect 10072 19008 10088 19072
rect 10152 19008 10160 19072
rect 9840 19007 10160 19008
rect 15770 19072 16090 19073
rect 15770 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15938 19072
rect 16002 19008 16018 19072
rect 16082 19008 16090 19072
rect 15770 19007 16090 19008
rect 6874 18528 7194 18529
rect 6874 18464 6882 18528
rect 6946 18464 6962 18528
rect 7026 18464 7042 18528
rect 7106 18464 7122 18528
rect 7186 18464 7194 18528
rect 6874 18463 7194 18464
rect 12805 18528 13125 18529
rect 12805 18464 12813 18528
rect 12877 18464 12893 18528
rect 12957 18464 12973 18528
rect 13037 18464 13053 18528
rect 13117 18464 13125 18528
rect 12805 18463 13125 18464
rect 3909 17984 4229 17985
rect 3909 17920 3917 17984
rect 3981 17920 3997 17984
rect 4061 17920 4077 17984
rect 4141 17920 4157 17984
rect 4221 17920 4229 17984
rect 3909 17919 4229 17920
rect 9840 17984 10160 17985
rect 9840 17920 9848 17984
rect 9912 17920 9928 17984
rect 9992 17920 10008 17984
rect 10072 17920 10088 17984
rect 10152 17920 10160 17984
rect 9840 17919 10160 17920
rect 15770 17984 16090 17985
rect 15770 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15938 17984
rect 16002 17920 16018 17984
rect 16082 17920 16090 17984
rect 15770 17919 16090 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 6874 17440 7194 17441
rect 6874 17376 6882 17440
rect 6946 17376 6962 17440
rect 7026 17376 7042 17440
rect 7106 17376 7122 17440
rect 7186 17376 7194 17440
rect 6874 17375 7194 17376
rect 12805 17440 13125 17441
rect 12805 17376 12813 17440
rect 12877 17376 12893 17440
rect 12957 17376 12973 17440
rect 13037 17376 13053 17440
rect 13117 17376 13125 17440
rect 12805 17375 13125 17376
rect 3909 16896 4229 16897
rect 3909 16832 3917 16896
rect 3981 16832 3997 16896
rect 4061 16832 4077 16896
rect 4141 16832 4157 16896
rect 4221 16832 4229 16896
rect 3909 16831 4229 16832
rect 9840 16896 10160 16897
rect 9840 16832 9848 16896
rect 9912 16832 9928 16896
rect 9992 16832 10008 16896
rect 10072 16832 10088 16896
rect 10152 16832 10160 16896
rect 9840 16831 10160 16832
rect 15770 16896 16090 16897
rect 15770 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15938 16896
rect 16002 16832 16018 16896
rect 16082 16832 16090 16896
rect 15770 16831 16090 16832
rect 6874 16352 7194 16353
rect 6874 16288 6882 16352
rect 6946 16288 6962 16352
rect 7026 16288 7042 16352
rect 7106 16288 7122 16352
rect 7186 16288 7194 16352
rect 6874 16287 7194 16288
rect 12805 16352 13125 16353
rect 12805 16288 12813 16352
rect 12877 16288 12893 16352
rect 12957 16288 12973 16352
rect 13037 16288 13053 16352
rect 13117 16288 13125 16352
rect 12805 16287 13125 16288
rect 3909 15808 4229 15809
rect 3909 15744 3917 15808
rect 3981 15744 3997 15808
rect 4061 15744 4077 15808
rect 4141 15744 4157 15808
rect 4221 15744 4229 15808
rect 3909 15743 4229 15744
rect 9840 15808 10160 15809
rect 9840 15744 9848 15808
rect 9912 15744 9928 15808
rect 9992 15744 10008 15808
rect 10072 15744 10088 15808
rect 10152 15744 10160 15808
rect 9840 15743 10160 15744
rect 15770 15808 16090 15809
rect 15770 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15938 15808
rect 16002 15744 16018 15808
rect 16082 15744 16090 15808
rect 15770 15743 16090 15744
rect 6085 15466 6151 15469
rect 7465 15466 7531 15469
rect 6085 15464 7531 15466
rect 6085 15408 6090 15464
rect 6146 15408 7470 15464
rect 7526 15408 7531 15464
rect 6085 15406 7531 15408
rect 6085 15403 6151 15406
rect 7465 15403 7531 15406
rect 6874 15264 7194 15265
rect 6874 15200 6882 15264
rect 6946 15200 6962 15264
rect 7026 15200 7042 15264
rect 7106 15200 7122 15264
rect 7186 15200 7194 15264
rect 6874 15199 7194 15200
rect 12805 15264 13125 15265
rect 12805 15200 12813 15264
rect 12877 15200 12893 15264
rect 12957 15200 12973 15264
rect 13037 15200 13053 15264
rect 13117 15200 13125 15264
rect 12805 15199 13125 15200
rect 3909 14720 4229 14721
rect 3909 14656 3917 14720
rect 3981 14656 3997 14720
rect 4061 14656 4077 14720
rect 4141 14656 4157 14720
rect 4221 14656 4229 14720
rect 3909 14655 4229 14656
rect 9840 14720 10160 14721
rect 9840 14656 9848 14720
rect 9912 14656 9928 14720
rect 9992 14656 10008 14720
rect 10072 14656 10088 14720
rect 10152 14656 10160 14720
rect 9840 14655 10160 14656
rect 15770 14720 16090 14721
rect 15770 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15938 14720
rect 16002 14656 16018 14720
rect 16082 14656 16090 14720
rect 15770 14655 16090 14656
rect 18137 14378 18203 14381
rect 19200 14378 20000 14408
rect 18137 14376 20000 14378
rect 18137 14320 18142 14376
rect 18198 14320 20000 14376
rect 18137 14318 20000 14320
rect 18137 14315 18203 14318
rect 19200 14288 20000 14318
rect 6874 14176 7194 14177
rect 6874 14112 6882 14176
rect 6946 14112 6962 14176
rect 7026 14112 7042 14176
rect 7106 14112 7122 14176
rect 7186 14112 7194 14176
rect 6874 14111 7194 14112
rect 12805 14176 13125 14177
rect 12805 14112 12813 14176
rect 12877 14112 12893 14176
rect 12957 14112 12973 14176
rect 13037 14112 13053 14176
rect 13117 14112 13125 14176
rect 12805 14111 13125 14112
rect 3909 13632 4229 13633
rect 3909 13568 3917 13632
rect 3981 13568 3997 13632
rect 4061 13568 4077 13632
rect 4141 13568 4157 13632
rect 4221 13568 4229 13632
rect 3909 13567 4229 13568
rect 9840 13632 10160 13633
rect 9840 13568 9848 13632
rect 9912 13568 9928 13632
rect 9992 13568 10008 13632
rect 10072 13568 10088 13632
rect 10152 13568 10160 13632
rect 9840 13567 10160 13568
rect 15770 13632 16090 13633
rect 15770 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15938 13632
rect 16002 13568 16018 13632
rect 16082 13568 16090 13632
rect 15770 13567 16090 13568
rect 6874 13088 7194 13089
rect 6874 13024 6882 13088
rect 6946 13024 6962 13088
rect 7026 13024 7042 13088
rect 7106 13024 7122 13088
rect 7186 13024 7194 13088
rect 6874 13023 7194 13024
rect 12805 13088 13125 13089
rect 12805 13024 12813 13088
rect 12877 13024 12893 13088
rect 12957 13024 12973 13088
rect 13037 13024 13053 13088
rect 13117 13024 13125 13088
rect 12805 13023 13125 13024
rect 3909 12544 4229 12545
rect 3909 12480 3917 12544
rect 3981 12480 3997 12544
rect 4061 12480 4077 12544
rect 4141 12480 4157 12544
rect 4221 12480 4229 12544
rect 3909 12479 4229 12480
rect 9840 12544 10160 12545
rect 9840 12480 9848 12544
rect 9912 12480 9928 12544
rect 9992 12480 10008 12544
rect 10072 12480 10088 12544
rect 10152 12480 10160 12544
rect 9840 12479 10160 12480
rect 15770 12544 16090 12545
rect 15770 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15938 12544
rect 16002 12480 16018 12544
rect 16082 12480 16090 12544
rect 15770 12479 16090 12480
rect 6874 12000 7194 12001
rect 6874 11936 6882 12000
rect 6946 11936 6962 12000
rect 7026 11936 7042 12000
rect 7106 11936 7122 12000
rect 7186 11936 7194 12000
rect 6874 11935 7194 11936
rect 12805 12000 13125 12001
rect 12805 11936 12813 12000
rect 12877 11936 12893 12000
rect 12957 11936 12973 12000
rect 13037 11936 13053 12000
rect 13117 11936 13125 12000
rect 12805 11935 13125 11936
rect 3909 11456 4229 11457
rect 3909 11392 3917 11456
rect 3981 11392 3997 11456
rect 4061 11392 4077 11456
rect 4141 11392 4157 11456
rect 4221 11392 4229 11456
rect 3909 11391 4229 11392
rect 9840 11456 10160 11457
rect 9840 11392 9848 11456
rect 9912 11392 9928 11456
rect 9992 11392 10008 11456
rect 10072 11392 10088 11456
rect 10152 11392 10160 11456
rect 9840 11391 10160 11392
rect 15770 11456 16090 11457
rect 15770 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15938 11456
rect 16002 11392 16018 11456
rect 16082 11392 16090 11456
rect 15770 11391 16090 11392
rect 6874 10912 7194 10913
rect 6874 10848 6882 10912
rect 6946 10848 6962 10912
rect 7026 10848 7042 10912
rect 7106 10848 7122 10912
rect 7186 10848 7194 10912
rect 6874 10847 7194 10848
rect 12805 10912 13125 10913
rect 12805 10848 12813 10912
rect 12877 10848 12893 10912
rect 12957 10848 12973 10912
rect 13037 10848 13053 10912
rect 13117 10848 13125 10912
rect 12805 10847 13125 10848
rect 3909 10368 4229 10369
rect 3909 10304 3917 10368
rect 3981 10304 3997 10368
rect 4061 10304 4077 10368
rect 4141 10304 4157 10368
rect 4221 10304 4229 10368
rect 3909 10303 4229 10304
rect 9840 10368 10160 10369
rect 9840 10304 9848 10368
rect 9912 10304 9928 10368
rect 9992 10304 10008 10368
rect 10072 10304 10088 10368
rect 10152 10304 10160 10368
rect 9840 10303 10160 10304
rect 15770 10368 16090 10369
rect 15770 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15938 10368
rect 16002 10304 16018 10368
rect 16082 10304 16090 10368
rect 15770 10303 16090 10304
rect 7005 10026 7071 10029
rect 8753 10026 8819 10029
rect 7005 10024 8819 10026
rect 7005 9968 7010 10024
rect 7066 9968 8758 10024
rect 8814 9968 8819 10024
rect 7005 9966 8819 9968
rect 7005 9963 7071 9966
rect 6874 9824 7194 9825
rect 6874 9760 6882 9824
rect 6946 9760 6962 9824
rect 7026 9760 7042 9824
rect 7106 9760 7122 9824
rect 7186 9760 7194 9824
rect 6874 9759 7194 9760
rect 7097 9690 7163 9693
rect 7422 9690 7482 9966
rect 8753 9963 8819 9966
rect 12805 9824 13125 9825
rect 12805 9760 12813 9824
rect 12877 9760 12893 9824
rect 12957 9760 12973 9824
rect 13037 9760 13053 9824
rect 13117 9760 13125 9824
rect 12805 9759 13125 9760
rect 7097 9688 7482 9690
rect 7097 9632 7102 9688
rect 7158 9632 7482 9688
rect 7097 9630 7482 9632
rect 7097 9627 7163 9630
rect 3909 9280 4229 9281
rect 3909 9216 3917 9280
rect 3981 9216 3997 9280
rect 4061 9216 4077 9280
rect 4141 9216 4157 9280
rect 4221 9216 4229 9280
rect 3909 9215 4229 9216
rect 9840 9280 10160 9281
rect 9840 9216 9848 9280
rect 9912 9216 9928 9280
rect 9992 9216 10008 9280
rect 10072 9216 10088 9280
rect 10152 9216 10160 9280
rect 9840 9215 10160 9216
rect 15770 9280 16090 9281
rect 15770 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15938 9280
rect 16002 9216 16018 9280
rect 16082 9216 16090 9280
rect 15770 9215 16090 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 6874 8736 7194 8737
rect 6874 8672 6882 8736
rect 6946 8672 6962 8736
rect 7026 8672 7042 8736
rect 7106 8672 7122 8736
rect 7186 8672 7194 8736
rect 6874 8671 7194 8672
rect 12805 8736 13125 8737
rect 12805 8672 12813 8736
rect 12877 8672 12893 8736
rect 12957 8672 12973 8736
rect 13037 8672 13053 8736
rect 13117 8672 13125 8736
rect 12805 8671 13125 8672
rect 3909 8192 4229 8193
rect 3909 8128 3917 8192
rect 3981 8128 3997 8192
rect 4061 8128 4077 8192
rect 4141 8128 4157 8192
rect 4221 8128 4229 8192
rect 3909 8127 4229 8128
rect 9840 8192 10160 8193
rect 9840 8128 9848 8192
rect 9912 8128 9928 8192
rect 9992 8128 10008 8192
rect 10072 8128 10088 8192
rect 10152 8128 10160 8192
rect 9840 8127 10160 8128
rect 15770 8192 16090 8193
rect 15770 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15938 8192
rect 16002 8128 16018 8192
rect 16082 8128 16090 8192
rect 15770 8127 16090 8128
rect 6874 7648 7194 7649
rect 6874 7584 6882 7648
rect 6946 7584 6962 7648
rect 7026 7584 7042 7648
rect 7106 7584 7122 7648
rect 7186 7584 7194 7648
rect 6874 7583 7194 7584
rect 12805 7648 13125 7649
rect 12805 7584 12813 7648
rect 12877 7584 12893 7648
rect 12957 7584 12973 7648
rect 13037 7584 13053 7648
rect 13117 7584 13125 7648
rect 12805 7583 13125 7584
rect 3909 7104 4229 7105
rect 3909 7040 3917 7104
rect 3981 7040 3997 7104
rect 4061 7040 4077 7104
rect 4141 7040 4157 7104
rect 4221 7040 4229 7104
rect 3909 7039 4229 7040
rect 9840 7104 10160 7105
rect 9840 7040 9848 7104
rect 9912 7040 9928 7104
rect 9992 7040 10008 7104
rect 10072 7040 10088 7104
rect 10152 7040 10160 7104
rect 9840 7039 10160 7040
rect 15770 7104 16090 7105
rect 15770 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15938 7104
rect 16002 7040 16018 7104
rect 16082 7040 16090 7104
rect 15770 7039 16090 7040
rect 6874 6560 7194 6561
rect 6874 6496 6882 6560
rect 6946 6496 6962 6560
rect 7026 6496 7042 6560
rect 7106 6496 7122 6560
rect 7186 6496 7194 6560
rect 6874 6495 7194 6496
rect 12805 6560 13125 6561
rect 12805 6496 12813 6560
rect 12877 6496 12893 6560
rect 12957 6496 12973 6560
rect 13037 6496 13053 6560
rect 13117 6496 13125 6560
rect 12805 6495 13125 6496
rect 3909 6016 4229 6017
rect 3909 5952 3917 6016
rect 3981 5952 3997 6016
rect 4061 5952 4077 6016
rect 4141 5952 4157 6016
rect 4221 5952 4229 6016
rect 3909 5951 4229 5952
rect 9840 6016 10160 6017
rect 9840 5952 9848 6016
rect 9912 5952 9928 6016
rect 9992 5952 10008 6016
rect 10072 5952 10088 6016
rect 10152 5952 10160 6016
rect 9840 5951 10160 5952
rect 15770 6016 16090 6017
rect 15770 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15938 6016
rect 16002 5952 16018 6016
rect 16082 5952 16090 6016
rect 15770 5951 16090 5952
rect 17861 5538 17927 5541
rect 19200 5538 20000 5568
rect 17861 5536 20000 5538
rect 17861 5480 17866 5536
rect 17922 5480 20000 5536
rect 17861 5478 20000 5480
rect 17861 5475 17927 5478
rect 6874 5472 7194 5473
rect 6874 5408 6882 5472
rect 6946 5408 6962 5472
rect 7026 5408 7042 5472
rect 7106 5408 7122 5472
rect 7186 5408 7194 5472
rect 6874 5407 7194 5408
rect 12805 5472 13125 5473
rect 12805 5408 12813 5472
rect 12877 5408 12893 5472
rect 12957 5408 12973 5472
rect 13037 5408 13053 5472
rect 13117 5408 13125 5472
rect 19200 5448 20000 5478
rect 12805 5407 13125 5408
rect 3909 4928 4229 4929
rect 3909 4864 3917 4928
rect 3981 4864 3997 4928
rect 4061 4864 4077 4928
rect 4141 4864 4157 4928
rect 4221 4864 4229 4928
rect 3909 4863 4229 4864
rect 9840 4928 10160 4929
rect 9840 4864 9848 4928
rect 9912 4864 9928 4928
rect 9992 4864 10008 4928
rect 10072 4864 10088 4928
rect 10152 4864 10160 4928
rect 9840 4863 10160 4864
rect 15770 4928 16090 4929
rect 15770 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15938 4928
rect 16002 4864 16018 4928
rect 16082 4864 16090 4928
rect 15770 4863 16090 4864
rect 6874 4384 7194 4385
rect 6874 4320 6882 4384
rect 6946 4320 6962 4384
rect 7026 4320 7042 4384
rect 7106 4320 7122 4384
rect 7186 4320 7194 4384
rect 6874 4319 7194 4320
rect 12805 4384 13125 4385
rect 12805 4320 12813 4384
rect 12877 4320 12893 4384
rect 12957 4320 12973 4384
rect 13037 4320 13053 4384
rect 13117 4320 13125 4384
rect 12805 4319 13125 4320
rect 3909 3840 4229 3841
rect 3909 3776 3917 3840
rect 3981 3776 3997 3840
rect 4061 3776 4077 3840
rect 4141 3776 4157 3840
rect 4221 3776 4229 3840
rect 3909 3775 4229 3776
rect 9840 3840 10160 3841
rect 9840 3776 9848 3840
rect 9912 3776 9928 3840
rect 9992 3776 10008 3840
rect 10072 3776 10088 3840
rect 10152 3776 10160 3840
rect 9840 3775 10160 3776
rect 15770 3840 16090 3841
rect 15770 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15938 3840
rect 16002 3776 16018 3840
rect 16082 3776 16090 3840
rect 15770 3775 16090 3776
rect 6874 3296 7194 3297
rect 6874 3232 6882 3296
rect 6946 3232 6962 3296
rect 7026 3232 7042 3296
rect 7106 3232 7122 3296
rect 7186 3232 7194 3296
rect 6874 3231 7194 3232
rect 12805 3296 13125 3297
rect 12805 3232 12813 3296
rect 12877 3232 12893 3296
rect 12957 3232 12973 3296
rect 13037 3232 13053 3296
rect 13117 3232 13125 3296
rect 12805 3231 13125 3232
rect 3909 2752 4229 2753
rect 3909 2688 3917 2752
rect 3981 2688 3997 2752
rect 4061 2688 4077 2752
rect 4141 2688 4157 2752
rect 4221 2688 4229 2752
rect 3909 2687 4229 2688
rect 9840 2752 10160 2753
rect 9840 2688 9848 2752
rect 9912 2688 9928 2752
rect 9992 2688 10008 2752
rect 10072 2688 10088 2752
rect 10152 2688 10160 2752
rect 9840 2687 10160 2688
rect 15770 2752 16090 2753
rect 15770 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15938 2752
rect 16002 2688 16018 2752
rect 16082 2688 16090 2752
rect 15770 2687 16090 2688
rect 6874 2208 7194 2209
rect 6874 2144 6882 2208
rect 6946 2144 6962 2208
rect 7026 2144 7042 2208
rect 7106 2144 7122 2208
rect 7186 2144 7194 2208
rect 6874 2143 7194 2144
rect 12805 2208 13125 2209
rect 12805 2144 12813 2208
rect 12877 2144 12893 2208
rect 12957 2144 12973 2208
rect 13037 2144 13053 2208
rect 13117 2144 13125 2208
rect 12805 2143 13125 2144
<< via3 >>
rect 3917 47356 3981 47360
rect 3917 47300 3921 47356
rect 3921 47300 3977 47356
rect 3977 47300 3981 47356
rect 3917 47296 3981 47300
rect 3997 47356 4061 47360
rect 3997 47300 4001 47356
rect 4001 47300 4057 47356
rect 4057 47300 4061 47356
rect 3997 47296 4061 47300
rect 4077 47356 4141 47360
rect 4077 47300 4081 47356
rect 4081 47300 4137 47356
rect 4137 47300 4141 47356
rect 4077 47296 4141 47300
rect 4157 47356 4221 47360
rect 4157 47300 4161 47356
rect 4161 47300 4217 47356
rect 4217 47300 4221 47356
rect 4157 47296 4221 47300
rect 9848 47356 9912 47360
rect 9848 47300 9852 47356
rect 9852 47300 9908 47356
rect 9908 47300 9912 47356
rect 9848 47296 9912 47300
rect 9928 47356 9992 47360
rect 9928 47300 9932 47356
rect 9932 47300 9988 47356
rect 9988 47300 9992 47356
rect 9928 47296 9992 47300
rect 10008 47356 10072 47360
rect 10008 47300 10012 47356
rect 10012 47300 10068 47356
rect 10068 47300 10072 47356
rect 10008 47296 10072 47300
rect 10088 47356 10152 47360
rect 10088 47300 10092 47356
rect 10092 47300 10148 47356
rect 10148 47300 10152 47356
rect 10088 47296 10152 47300
rect 15778 47356 15842 47360
rect 15778 47300 15782 47356
rect 15782 47300 15838 47356
rect 15838 47300 15842 47356
rect 15778 47296 15842 47300
rect 15858 47356 15922 47360
rect 15858 47300 15862 47356
rect 15862 47300 15918 47356
rect 15918 47300 15922 47356
rect 15858 47296 15922 47300
rect 15938 47356 16002 47360
rect 15938 47300 15942 47356
rect 15942 47300 15998 47356
rect 15998 47300 16002 47356
rect 15938 47296 16002 47300
rect 16018 47356 16082 47360
rect 16018 47300 16022 47356
rect 16022 47300 16078 47356
rect 16078 47300 16082 47356
rect 16018 47296 16082 47300
rect 6882 46812 6946 46816
rect 6882 46756 6886 46812
rect 6886 46756 6942 46812
rect 6942 46756 6946 46812
rect 6882 46752 6946 46756
rect 6962 46812 7026 46816
rect 6962 46756 6966 46812
rect 6966 46756 7022 46812
rect 7022 46756 7026 46812
rect 6962 46752 7026 46756
rect 7042 46812 7106 46816
rect 7042 46756 7046 46812
rect 7046 46756 7102 46812
rect 7102 46756 7106 46812
rect 7042 46752 7106 46756
rect 7122 46812 7186 46816
rect 7122 46756 7126 46812
rect 7126 46756 7182 46812
rect 7182 46756 7186 46812
rect 7122 46752 7186 46756
rect 12813 46812 12877 46816
rect 12813 46756 12817 46812
rect 12817 46756 12873 46812
rect 12873 46756 12877 46812
rect 12813 46752 12877 46756
rect 12893 46812 12957 46816
rect 12893 46756 12897 46812
rect 12897 46756 12953 46812
rect 12953 46756 12957 46812
rect 12893 46752 12957 46756
rect 12973 46812 13037 46816
rect 12973 46756 12977 46812
rect 12977 46756 13033 46812
rect 13033 46756 13037 46812
rect 12973 46752 13037 46756
rect 13053 46812 13117 46816
rect 13053 46756 13057 46812
rect 13057 46756 13113 46812
rect 13113 46756 13117 46812
rect 13053 46752 13117 46756
rect 3917 46268 3981 46272
rect 3917 46212 3921 46268
rect 3921 46212 3977 46268
rect 3977 46212 3981 46268
rect 3917 46208 3981 46212
rect 3997 46268 4061 46272
rect 3997 46212 4001 46268
rect 4001 46212 4057 46268
rect 4057 46212 4061 46268
rect 3997 46208 4061 46212
rect 4077 46268 4141 46272
rect 4077 46212 4081 46268
rect 4081 46212 4137 46268
rect 4137 46212 4141 46268
rect 4077 46208 4141 46212
rect 4157 46268 4221 46272
rect 4157 46212 4161 46268
rect 4161 46212 4217 46268
rect 4217 46212 4221 46268
rect 4157 46208 4221 46212
rect 9848 46268 9912 46272
rect 9848 46212 9852 46268
rect 9852 46212 9908 46268
rect 9908 46212 9912 46268
rect 9848 46208 9912 46212
rect 9928 46268 9992 46272
rect 9928 46212 9932 46268
rect 9932 46212 9988 46268
rect 9988 46212 9992 46268
rect 9928 46208 9992 46212
rect 10008 46268 10072 46272
rect 10008 46212 10012 46268
rect 10012 46212 10068 46268
rect 10068 46212 10072 46268
rect 10008 46208 10072 46212
rect 10088 46268 10152 46272
rect 10088 46212 10092 46268
rect 10092 46212 10148 46268
rect 10148 46212 10152 46268
rect 10088 46208 10152 46212
rect 15778 46268 15842 46272
rect 15778 46212 15782 46268
rect 15782 46212 15838 46268
rect 15838 46212 15842 46268
rect 15778 46208 15842 46212
rect 15858 46268 15922 46272
rect 15858 46212 15862 46268
rect 15862 46212 15918 46268
rect 15918 46212 15922 46268
rect 15858 46208 15922 46212
rect 15938 46268 16002 46272
rect 15938 46212 15942 46268
rect 15942 46212 15998 46268
rect 15998 46212 16002 46268
rect 15938 46208 16002 46212
rect 16018 46268 16082 46272
rect 16018 46212 16022 46268
rect 16022 46212 16078 46268
rect 16078 46212 16082 46268
rect 16018 46208 16082 46212
rect 6882 45724 6946 45728
rect 6882 45668 6886 45724
rect 6886 45668 6942 45724
rect 6942 45668 6946 45724
rect 6882 45664 6946 45668
rect 6962 45724 7026 45728
rect 6962 45668 6966 45724
rect 6966 45668 7022 45724
rect 7022 45668 7026 45724
rect 6962 45664 7026 45668
rect 7042 45724 7106 45728
rect 7042 45668 7046 45724
rect 7046 45668 7102 45724
rect 7102 45668 7106 45724
rect 7042 45664 7106 45668
rect 7122 45724 7186 45728
rect 7122 45668 7126 45724
rect 7126 45668 7182 45724
rect 7182 45668 7186 45724
rect 7122 45664 7186 45668
rect 12813 45724 12877 45728
rect 12813 45668 12817 45724
rect 12817 45668 12873 45724
rect 12873 45668 12877 45724
rect 12813 45664 12877 45668
rect 12893 45724 12957 45728
rect 12893 45668 12897 45724
rect 12897 45668 12953 45724
rect 12953 45668 12957 45724
rect 12893 45664 12957 45668
rect 12973 45724 13037 45728
rect 12973 45668 12977 45724
rect 12977 45668 13033 45724
rect 13033 45668 13037 45724
rect 12973 45664 13037 45668
rect 13053 45724 13117 45728
rect 13053 45668 13057 45724
rect 13057 45668 13113 45724
rect 13113 45668 13117 45724
rect 13053 45664 13117 45668
rect 3917 45180 3981 45184
rect 3917 45124 3921 45180
rect 3921 45124 3977 45180
rect 3977 45124 3981 45180
rect 3917 45120 3981 45124
rect 3997 45180 4061 45184
rect 3997 45124 4001 45180
rect 4001 45124 4057 45180
rect 4057 45124 4061 45180
rect 3997 45120 4061 45124
rect 4077 45180 4141 45184
rect 4077 45124 4081 45180
rect 4081 45124 4137 45180
rect 4137 45124 4141 45180
rect 4077 45120 4141 45124
rect 4157 45180 4221 45184
rect 4157 45124 4161 45180
rect 4161 45124 4217 45180
rect 4217 45124 4221 45180
rect 4157 45120 4221 45124
rect 9848 45180 9912 45184
rect 9848 45124 9852 45180
rect 9852 45124 9908 45180
rect 9908 45124 9912 45180
rect 9848 45120 9912 45124
rect 9928 45180 9992 45184
rect 9928 45124 9932 45180
rect 9932 45124 9988 45180
rect 9988 45124 9992 45180
rect 9928 45120 9992 45124
rect 10008 45180 10072 45184
rect 10008 45124 10012 45180
rect 10012 45124 10068 45180
rect 10068 45124 10072 45180
rect 10008 45120 10072 45124
rect 10088 45180 10152 45184
rect 10088 45124 10092 45180
rect 10092 45124 10148 45180
rect 10148 45124 10152 45180
rect 10088 45120 10152 45124
rect 15778 45180 15842 45184
rect 15778 45124 15782 45180
rect 15782 45124 15838 45180
rect 15838 45124 15842 45180
rect 15778 45120 15842 45124
rect 15858 45180 15922 45184
rect 15858 45124 15862 45180
rect 15862 45124 15918 45180
rect 15918 45124 15922 45180
rect 15858 45120 15922 45124
rect 15938 45180 16002 45184
rect 15938 45124 15942 45180
rect 15942 45124 15998 45180
rect 15998 45124 16002 45180
rect 15938 45120 16002 45124
rect 16018 45180 16082 45184
rect 16018 45124 16022 45180
rect 16022 45124 16078 45180
rect 16078 45124 16082 45180
rect 16018 45120 16082 45124
rect 6882 44636 6946 44640
rect 6882 44580 6886 44636
rect 6886 44580 6942 44636
rect 6942 44580 6946 44636
rect 6882 44576 6946 44580
rect 6962 44636 7026 44640
rect 6962 44580 6966 44636
rect 6966 44580 7022 44636
rect 7022 44580 7026 44636
rect 6962 44576 7026 44580
rect 7042 44636 7106 44640
rect 7042 44580 7046 44636
rect 7046 44580 7102 44636
rect 7102 44580 7106 44636
rect 7042 44576 7106 44580
rect 7122 44636 7186 44640
rect 7122 44580 7126 44636
rect 7126 44580 7182 44636
rect 7182 44580 7186 44636
rect 7122 44576 7186 44580
rect 12813 44636 12877 44640
rect 12813 44580 12817 44636
rect 12817 44580 12873 44636
rect 12873 44580 12877 44636
rect 12813 44576 12877 44580
rect 12893 44636 12957 44640
rect 12893 44580 12897 44636
rect 12897 44580 12953 44636
rect 12953 44580 12957 44636
rect 12893 44576 12957 44580
rect 12973 44636 13037 44640
rect 12973 44580 12977 44636
rect 12977 44580 13033 44636
rect 13033 44580 13037 44636
rect 12973 44576 13037 44580
rect 13053 44636 13117 44640
rect 13053 44580 13057 44636
rect 13057 44580 13113 44636
rect 13113 44580 13117 44636
rect 13053 44576 13117 44580
rect 3917 44092 3981 44096
rect 3917 44036 3921 44092
rect 3921 44036 3977 44092
rect 3977 44036 3981 44092
rect 3917 44032 3981 44036
rect 3997 44092 4061 44096
rect 3997 44036 4001 44092
rect 4001 44036 4057 44092
rect 4057 44036 4061 44092
rect 3997 44032 4061 44036
rect 4077 44092 4141 44096
rect 4077 44036 4081 44092
rect 4081 44036 4137 44092
rect 4137 44036 4141 44092
rect 4077 44032 4141 44036
rect 4157 44092 4221 44096
rect 4157 44036 4161 44092
rect 4161 44036 4217 44092
rect 4217 44036 4221 44092
rect 4157 44032 4221 44036
rect 9848 44092 9912 44096
rect 9848 44036 9852 44092
rect 9852 44036 9908 44092
rect 9908 44036 9912 44092
rect 9848 44032 9912 44036
rect 9928 44092 9992 44096
rect 9928 44036 9932 44092
rect 9932 44036 9988 44092
rect 9988 44036 9992 44092
rect 9928 44032 9992 44036
rect 10008 44092 10072 44096
rect 10008 44036 10012 44092
rect 10012 44036 10068 44092
rect 10068 44036 10072 44092
rect 10008 44032 10072 44036
rect 10088 44092 10152 44096
rect 10088 44036 10092 44092
rect 10092 44036 10148 44092
rect 10148 44036 10152 44092
rect 10088 44032 10152 44036
rect 15778 44092 15842 44096
rect 15778 44036 15782 44092
rect 15782 44036 15838 44092
rect 15838 44036 15842 44092
rect 15778 44032 15842 44036
rect 15858 44092 15922 44096
rect 15858 44036 15862 44092
rect 15862 44036 15918 44092
rect 15918 44036 15922 44092
rect 15858 44032 15922 44036
rect 15938 44092 16002 44096
rect 15938 44036 15942 44092
rect 15942 44036 15998 44092
rect 15998 44036 16002 44092
rect 15938 44032 16002 44036
rect 16018 44092 16082 44096
rect 16018 44036 16022 44092
rect 16022 44036 16078 44092
rect 16078 44036 16082 44092
rect 16018 44032 16082 44036
rect 6882 43548 6946 43552
rect 6882 43492 6886 43548
rect 6886 43492 6942 43548
rect 6942 43492 6946 43548
rect 6882 43488 6946 43492
rect 6962 43548 7026 43552
rect 6962 43492 6966 43548
rect 6966 43492 7022 43548
rect 7022 43492 7026 43548
rect 6962 43488 7026 43492
rect 7042 43548 7106 43552
rect 7042 43492 7046 43548
rect 7046 43492 7102 43548
rect 7102 43492 7106 43548
rect 7042 43488 7106 43492
rect 7122 43548 7186 43552
rect 7122 43492 7126 43548
rect 7126 43492 7182 43548
rect 7182 43492 7186 43548
rect 7122 43488 7186 43492
rect 12813 43548 12877 43552
rect 12813 43492 12817 43548
rect 12817 43492 12873 43548
rect 12873 43492 12877 43548
rect 12813 43488 12877 43492
rect 12893 43548 12957 43552
rect 12893 43492 12897 43548
rect 12897 43492 12953 43548
rect 12953 43492 12957 43548
rect 12893 43488 12957 43492
rect 12973 43548 13037 43552
rect 12973 43492 12977 43548
rect 12977 43492 13033 43548
rect 13033 43492 13037 43548
rect 12973 43488 13037 43492
rect 13053 43548 13117 43552
rect 13053 43492 13057 43548
rect 13057 43492 13113 43548
rect 13113 43492 13117 43548
rect 13053 43488 13117 43492
rect 3917 43004 3981 43008
rect 3917 42948 3921 43004
rect 3921 42948 3977 43004
rect 3977 42948 3981 43004
rect 3917 42944 3981 42948
rect 3997 43004 4061 43008
rect 3997 42948 4001 43004
rect 4001 42948 4057 43004
rect 4057 42948 4061 43004
rect 3997 42944 4061 42948
rect 4077 43004 4141 43008
rect 4077 42948 4081 43004
rect 4081 42948 4137 43004
rect 4137 42948 4141 43004
rect 4077 42944 4141 42948
rect 4157 43004 4221 43008
rect 4157 42948 4161 43004
rect 4161 42948 4217 43004
rect 4217 42948 4221 43004
rect 4157 42944 4221 42948
rect 9848 43004 9912 43008
rect 9848 42948 9852 43004
rect 9852 42948 9908 43004
rect 9908 42948 9912 43004
rect 9848 42944 9912 42948
rect 9928 43004 9992 43008
rect 9928 42948 9932 43004
rect 9932 42948 9988 43004
rect 9988 42948 9992 43004
rect 9928 42944 9992 42948
rect 10008 43004 10072 43008
rect 10008 42948 10012 43004
rect 10012 42948 10068 43004
rect 10068 42948 10072 43004
rect 10008 42944 10072 42948
rect 10088 43004 10152 43008
rect 10088 42948 10092 43004
rect 10092 42948 10148 43004
rect 10148 42948 10152 43004
rect 10088 42944 10152 42948
rect 15778 43004 15842 43008
rect 15778 42948 15782 43004
rect 15782 42948 15838 43004
rect 15838 42948 15842 43004
rect 15778 42944 15842 42948
rect 15858 43004 15922 43008
rect 15858 42948 15862 43004
rect 15862 42948 15918 43004
rect 15918 42948 15922 43004
rect 15858 42944 15922 42948
rect 15938 43004 16002 43008
rect 15938 42948 15942 43004
rect 15942 42948 15998 43004
rect 15998 42948 16002 43004
rect 15938 42944 16002 42948
rect 16018 43004 16082 43008
rect 16018 42948 16022 43004
rect 16022 42948 16078 43004
rect 16078 42948 16082 43004
rect 16018 42944 16082 42948
rect 6882 42460 6946 42464
rect 6882 42404 6886 42460
rect 6886 42404 6942 42460
rect 6942 42404 6946 42460
rect 6882 42400 6946 42404
rect 6962 42460 7026 42464
rect 6962 42404 6966 42460
rect 6966 42404 7022 42460
rect 7022 42404 7026 42460
rect 6962 42400 7026 42404
rect 7042 42460 7106 42464
rect 7042 42404 7046 42460
rect 7046 42404 7102 42460
rect 7102 42404 7106 42460
rect 7042 42400 7106 42404
rect 7122 42460 7186 42464
rect 7122 42404 7126 42460
rect 7126 42404 7182 42460
rect 7182 42404 7186 42460
rect 7122 42400 7186 42404
rect 12813 42460 12877 42464
rect 12813 42404 12817 42460
rect 12817 42404 12873 42460
rect 12873 42404 12877 42460
rect 12813 42400 12877 42404
rect 12893 42460 12957 42464
rect 12893 42404 12897 42460
rect 12897 42404 12953 42460
rect 12953 42404 12957 42460
rect 12893 42400 12957 42404
rect 12973 42460 13037 42464
rect 12973 42404 12977 42460
rect 12977 42404 13033 42460
rect 13033 42404 13037 42460
rect 12973 42400 13037 42404
rect 13053 42460 13117 42464
rect 13053 42404 13057 42460
rect 13057 42404 13113 42460
rect 13113 42404 13117 42460
rect 13053 42400 13117 42404
rect 3917 41916 3981 41920
rect 3917 41860 3921 41916
rect 3921 41860 3977 41916
rect 3977 41860 3981 41916
rect 3917 41856 3981 41860
rect 3997 41916 4061 41920
rect 3997 41860 4001 41916
rect 4001 41860 4057 41916
rect 4057 41860 4061 41916
rect 3997 41856 4061 41860
rect 4077 41916 4141 41920
rect 4077 41860 4081 41916
rect 4081 41860 4137 41916
rect 4137 41860 4141 41916
rect 4077 41856 4141 41860
rect 4157 41916 4221 41920
rect 4157 41860 4161 41916
rect 4161 41860 4217 41916
rect 4217 41860 4221 41916
rect 4157 41856 4221 41860
rect 9848 41916 9912 41920
rect 9848 41860 9852 41916
rect 9852 41860 9908 41916
rect 9908 41860 9912 41916
rect 9848 41856 9912 41860
rect 9928 41916 9992 41920
rect 9928 41860 9932 41916
rect 9932 41860 9988 41916
rect 9988 41860 9992 41916
rect 9928 41856 9992 41860
rect 10008 41916 10072 41920
rect 10008 41860 10012 41916
rect 10012 41860 10068 41916
rect 10068 41860 10072 41916
rect 10008 41856 10072 41860
rect 10088 41916 10152 41920
rect 10088 41860 10092 41916
rect 10092 41860 10148 41916
rect 10148 41860 10152 41916
rect 10088 41856 10152 41860
rect 15778 41916 15842 41920
rect 15778 41860 15782 41916
rect 15782 41860 15838 41916
rect 15838 41860 15842 41916
rect 15778 41856 15842 41860
rect 15858 41916 15922 41920
rect 15858 41860 15862 41916
rect 15862 41860 15918 41916
rect 15918 41860 15922 41916
rect 15858 41856 15922 41860
rect 15938 41916 16002 41920
rect 15938 41860 15942 41916
rect 15942 41860 15998 41916
rect 15998 41860 16002 41916
rect 15938 41856 16002 41860
rect 16018 41916 16082 41920
rect 16018 41860 16022 41916
rect 16022 41860 16078 41916
rect 16078 41860 16082 41916
rect 16018 41856 16082 41860
rect 6882 41372 6946 41376
rect 6882 41316 6886 41372
rect 6886 41316 6942 41372
rect 6942 41316 6946 41372
rect 6882 41312 6946 41316
rect 6962 41372 7026 41376
rect 6962 41316 6966 41372
rect 6966 41316 7022 41372
rect 7022 41316 7026 41372
rect 6962 41312 7026 41316
rect 7042 41372 7106 41376
rect 7042 41316 7046 41372
rect 7046 41316 7102 41372
rect 7102 41316 7106 41372
rect 7042 41312 7106 41316
rect 7122 41372 7186 41376
rect 7122 41316 7126 41372
rect 7126 41316 7182 41372
rect 7182 41316 7186 41372
rect 7122 41312 7186 41316
rect 12813 41372 12877 41376
rect 12813 41316 12817 41372
rect 12817 41316 12873 41372
rect 12873 41316 12877 41372
rect 12813 41312 12877 41316
rect 12893 41372 12957 41376
rect 12893 41316 12897 41372
rect 12897 41316 12953 41372
rect 12953 41316 12957 41372
rect 12893 41312 12957 41316
rect 12973 41372 13037 41376
rect 12973 41316 12977 41372
rect 12977 41316 13033 41372
rect 13033 41316 13037 41372
rect 12973 41312 13037 41316
rect 13053 41372 13117 41376
rect 13053 41316 13057 41372
rect 13057 41316 13113 41372
rect 13113 41316 13117 41372
rect 13053 41312 13117 41316
rect 3917 40828 3981 40832
rect 3917 40772 3921 40828
rect 3921 40772 3977 40828
rect 3977 40772 3981 40828
rect 3917 40768 3981 40772
rect 3997 40828 4061 40832
rect 3997 40772 4001 40828
rect 4001 40772 4057 40828
rect 4057 40772 4061 40828
rect 3997 40768 4061 40772
rect 4077 40828 4141 40832
rect 4077 40772 4081 40828
rect 4081 40772 4137 40828
rect 4137 40772 4141 40828
rect 4077 40768 4141 40772
rect 4157 40828 4221 40832
rect 4157 40772 4161 40828
rect 4161 40772 4217 40828
rect 4217 40772 4221 40828
rect 4157 40768 4221 40772
rect 9848 40828 9912 40832
rect 9848 40772 9852 40828
rect 9852 40772 9908 40828
rect 9908 40772 9912 40828
rect 9848 40768 9912 40772
rect 9928 40828 9992 40832
rect 9928 40772 9932 40828
rect 9932 40772 9988 40828
rect 9988 40772 9992 40828
rect 9928 40768 9992 40772
rect 10008 40828 10072 40832
rect 10008 40772 10012 40828
rect 10012 40772 10068 40828
rect 10068 40772 10072 40828
rect 10008 40768 10072 40772
rect 10088 40828 10152 40832
rect 10088 40772 10092 40828
rect 10092 40772 10148 40828
rect 10148 40772 10152 40828
rect 10088 40768 10152 40772
rect 15778 40828 15842 40832
rect 15778 40772 15782 40828
rect 15782 40772 15838 40828
rect 15838 40772 15842 40828
rect 15778 40768 15842 40772
rect 15858 40828 15922 40832
rect 15858 40772 15862 40828
rect 15862 40772 15918 40828
rect 15918 40772 15922 40828
rect 15858 40768 15922 40772
rect 15938 40828 16002 40832
rect 15938 40772 15942 40828
rect 15942 40772 15998 40828
rect 15998 40772 16002 40828
rect 15938 40768 16002 40772
rect 16018 40828 16082 40832
rect 16018 40772 16022 40828
rect 16022 40772 16078 40828
rect 16078 40772 16082 40828
rect 16018 40768 16082 40772
rect 6882 40284 6946 40288
rect 6882 40228 6886 40284
rect 6886 40228 6942 40284
rect 6942 40228 6946 40284
rect 6882 40224 6946 40228
rect 6962 40284 7026 40288
rect 6962 40228 6966 40284
rect 6966 40228 7022 40284
rect 7022 40228 7026 40284
rect 6962 40224 7026 40228
rect 7042 40284 7106 40288
rect 7042 40228 7046 40284
rect 7046 40228 7102 40284
rect 7102 40228 7106 40284
rect 7042 40224 7106 40228
rect 7122 40284 7186 40288
rect 7122 40228 7126 40284
rect 7126 40228 7182 40284
rect 7182 40228 7186 40284
rect 7122 40224 7186 40228
rect 12813 40284 12877 40288
rect 12813 40228 12817 40284
rect 12817 40228 12873 40284
rect 12873 40228 12877 40284
rect 12813 40224 12877 40228
rect 12893 40284 12957 40288
rect 12893 40228 12897 40284
rect 12897 40228 12953 40284
rect 12953 40228 12957 40284
rect 12893 40224 12957 40228
rect 12973 40284 13037 40288
rect 12973 40228 12977 40284
rect 12977 40228 13033 40284
rect 13033 40228 13037 40284
rect 12973 40224 13037 40228
rect 13053 40284 13117 40288
rect 13053 40228 13057 40284
rect 13057 40228 13113 40284
rect 13113 40228 13117 40284
rect 13053 40224 13117 40228
rect 3917 39740 3981 39744
rect 3917 39684 3921 39740
rect 3921 39684 3977 39740
rect 3977 39684 3981 39740
rect 3917 39680 3981 39684
rect 3997 39740 4061 39744
rect 3997 39684 4001 39740
rect 4001 39684 4057 39740
rect 4057 39684 4061 39740
rect 3997 39680 4061 39684
rect 4077 39740 4141 39744
rect 4077 39684 4081 39740
rect 4081 39684 4137 39740
rect 4137 39684 4141 39740
rect 4077 39680 4141 39684
rect 4157 39740 4221 39744
rect 4157 39684 4161 39740
rect 4161 39684 4217 39740
rect 4217 39684 4221 39740
rect 4157 39680 4221 39684
rect 9848 39740 9912 39744
rect 9848 39684 9852 39740
rect 9852 39684 9908 39740
rect 9908 39684 9912 39740
rect 9848 39680 9912 39684
rect 9928 39740 9992 39744
rect 9928 39684 9932 39740
rect 9932 39684 9988 39740
rect 9988 39684 9992 39740
rect 9928 39680 9992 39684
rect 10008 39740 10072 39744
rect 10008 39684 10012 39740
rect 10012 39684 10068 39740
rect 10068 39684 10072 39740
rect 10008 39680 10072 39684
rect 10088 39740 10152 39744
rect 10088 39684 10092 39740
rect 10092 39684 10148 39740
rect 10148 39684 10152 39740
rect 10088 39680 10152 39684
rect 15778 39740 15842 39744
rect 15778 39684 15782 39740
rect 15782 39684 15838 39740
rect 15838 39684 15842 39740
rect 15778 39680 15842 39684
rect 15858 39740 15922 39744
rect 15858 39684 15862 39740
rect 15862 39684 15918 39740
rect 15918 39684 15922 39740
rect 15858 39680 15922 39684
rect 15938 39740 16002 39744
rect 15938 39684 15942 39740
rect 15942 39684 15998 39740
rect 15998 39684 16002 39740
rect 15938 39680 16002 39684
rect 16018 39740 16082 39744
rect 16018 39684 16022 39740
rect 16022 39684 16078 39740
rect 16078 39684 16082 39740
rect 16018 39680 16082 39684
rect 6882 39196 6946 39200
rect 6882 39140 6886 39196
rect 6886 39140 6942 39196
rect 6942 39140 6946 39196
rect 6882 39136 6946 39140
rect 6962 39196 7026 39200
rect 6962 39140 6966 39196
rect 6966 39140 7022 39196
rect 7022 39140 7026 39196
rect 6962 39136 7026 39140
rect 7042 39196 7106 39200
rect 7042 39140 7046 39196
rect 7046 39140 7102 39196
rect 7102 39140 7106 39196
rect 7042 39136 7106 39140
rect 7122 39196 7186 39200
rect 7122 39140 7126 39196
rect 7126 39140 7182 39196
rect 7182 39140 7186 39196
rect 7122 39136 7186 39140
rect 12813 39196 12877 39200
rect 12813 39140 12817 39196
rect 12817 39140 12873 39196
rect 12873 39140 12877 39196
rect 12813 39136 12877 39140
rect 12893 39196 12957 39200
rect 12893 39140 12897 39196
rect 12897 39140 12953 39196
rect 12953 39140 12957 39196
rect 12893 39136 12957 39140
rect 12973 39196 13037 39200
rect 12973 39140 12977 39196
rect 12977 39140 13033 39196
rect 13033 39140 13037 39196
rect 12973 39136 13037 39140
rect 13053 39196 13117 39200
rect 13053 39140 13057 39196
rect 13057 39140 13113 39196
rect 13113 39140 13117 39196
rect 13053 39136 13117 39140
rect 3917 38652 3981 38656
rect 3917 38596 3921 38652
rect 3921 38596 3977 38652
rect 3977 38596 3981 38652
rect 3917 38592 3981 38596
rect 3997 38652 4061 38656
rect 3997 38596 4001 38652
rect 4001 38596 4057 38652
rect 4057 38596 4061 38652
rect 3997 38592 4061 38596
rect 4077 38652 4141 38656
rect 4077 38596 4081 38652
rect 4081 38596 4137 38652
rect 4137 38596 4141 38652
rect 4077 38592 4141 38596
rect 4157 38652 4221 38656
rect 4157 38596 4161 38652
rect 4161 38596 4217 38652
rect 4217 38596 4221 38652
rect 4157 38592 4221 38596
rect 9848 38652 9912 38656
rect 9848 38596 9852 38652
rect 9852 38596 9908 38652
rect 9908 38596 9912 38652
rect 9848 38592 9912 38596
rect 9928 38652 9992 38656
rect 9928 38596 9932 38652
rect 9932 38596 9988 38652
rect 9988 38596 9992 38652
rect 9928 38592 9992 38596
rect 10008 38652 10072 38656
rect 10008 38596 10012 38652
rect 10012 38596 10068 38652
rect 10068 38596 10072 38652
rect 10008 38592 10072 38596
rect 10088 38652 10152 38656
rect 10088 38596 10092 38652
rect 10092 38596 10148 38652
rect 10148 38596 10152 38652
rect 10088 38592 10152 38596
rect 15778 38652 15842 38656
rect 15778 38596 15782 38652
rect 15782 38596 15838 38652
rect 15838 38596 15842 38652
rect 15778 38592 15842 38596
rect 15858 38652 15922 38656
rect 15858 38596 15862 38652
rect 15862 38596 15918 38652
rect 15918 38596 15922 38652
rect 15858 38592 15922 38596
rect 15938 38652 16002 38656
rect 15938 38596 15942 38652
rect 15942 38596 15998 38652
rect 15998 38596 16002 38652
rect 15938 38592 16002 38596
rect 16018 38652 16082 38656
rect 16018 38596 16022 38652
rect 16022 38596 16078 38652
rect 16078 38596 16082 38652
rect 16018 38592 16082 38596
rect 6882 38108 6946 38112
rect 6882 38052 6886 38108
rect 6886 38052 6942 38108
rect 6942 38052 6946 38108
rect 6882 38048 6946 38052
rect 6962 38108 7026 38112
rect 6962 38052 6966 38108
rect 6966 38052 7022 38108
rect 7022 38052 7026 38108
rect 6962 38048 7026 38052
rect 7042 38108 7106 38112
rect 7042 38052 7046 38108
rect 7046 38052 7102 38108
rect 7102 38052 7106 38108
rect 7042 38048 7106 38052
rect 7122 38108 7186 38112
rect 7122 38052 7126 38108
rect 7126 38052 7182 38108
rect 7182 38052 7186 38108
rect 7122 38048 7186 38052
rect 12813 38108 12877 38112
rect 12813 38052 12817 38108
rect 12817 38052 12873 38108
rect 12873 38052 12877 38108
rect 12813 38048 12877 38052
rect 12893 38108 12957 38112
rect 12893 38052 12897 38108
rect 12897 38052 12953 38108
rect 12953 38052 12957 38108
rect 12893 38048 12957 38052
rect 12973 38108 13037 38112
rect 12973 38052 12977 38108
rect 12977 38052 13033 38108
rect 13033 38052 13037 38108
rect 12973 38048 13037 38052
rect 13053 38108 13117 38112
rect 13053 38052 13057 38108
rect 13057 38052 13113 38108
rect 13113 38052 13117 38108
rect 13053 38048 13117 38052
rect 3917 37564 3981 37568
rect 3917 37508 3921 37564
rect 3921 37508 3977 37564
rect 3977 37508 3981 37564
rect 3917 37504 3981 37508
rect 3997 37564 4061 37568
rect 3997 37508 4001 37564
rect 4001 37508 4057 37564
rect 4057 37508 4061 37564
rect 3997 37504 4061 37508
rect 4077 37564 4141 37568
rect 4077 37508 4081 37564
rect 4081 37508 4137 37564
rect 4137 37508 4141 37564
rect 4077 37504 4141 37508
rect 4157 37564 4221 37568
rect 4157 37508 4161 37564
rect 4161 37508 4217 37564
rect 4217 37508 4221 37564
rect 4157 37504 4221 37508
rect 9848 37564 9912 37568
rect 9848 37508 9852 37564
rect 9852 37508 9908 37564
rect 9908 37508 9912 37564
rect 9848 37504 9912 37508
rect 9928 37564 9992 37568
rect 9928 37508 9932 37564
rect 9932 37508 9988 37564
rect 9988 37508 9992 37564
rect 9928 37504 9992 37508
rect 10008 37564 10072 37568
rect 10008 37508 10012 37564
rect 10012 37508 10068 37564
rect 10068 37508 10072 37564
rect 10008 37504 10072 37508
rect 10088 37564 10152 37568
rect 10088 37508 10092 37564
rect 10092 37508 10148 37564
rect 10148 37508 10152 37564
rect 10088 37504 10152 37508
rect 15778 37564 15842 37568
rect 15778 37508 15782 37564
rect 15782 37508 15838 37564
rect 15838 37508 15842 37564
rect 15778 37504 15842 37508
rect 15858 37564 15922 37568
rect 15858 37508 15862 37564
rect 15862 37508 15918 37564
rect 15918 37508 15922 37564
rect 15858 37504 15922 37508
rect 15938 37564 16002 37568
rect 15938 37508 15942 37564
rect 15942 37508 15998 37564
rect 15998 37508 16002 37564
rect 15938 37504 16002 37508
rect 16018 37564 16082 37568
rect 16018 37508 16022 37564
rect 16022 37508 16078 37564
rect 16078 37508 16082 37564
rect 16018 37504 16082 37508
rect 6882 37020 6946 37024
rect 6882 36964 6886 37020
rect 6886 36964 6942 37020
rect 6942 36964 6946 37020
rect 6882 36960 6946 36964
rect 6962 37020 7026 37024
rect 6962 36964 6966 37020
rect 6966 36964 7022 37020
rect 7022 36964 7026 37020
rect 6962 36960 7026 36964
rect 7042 37020 7106 37024
rect 7042 36964 7046 37020
rect 7046 36964 7102 37020
rect 7102 36964 7106 37020
rect 7042 36960 7106 36964
rect 7122 37020 7186 37024
rect 7122 36964 7126 37020
rect 7126 36964 7182 37020
rect 7182 36964 7186 37020
rect 7122 36960 7186 36964
rect 12813 37020 12877 37024
rect 12813 36964 12817 37020
rect 12817 36964 12873 37020
rect 12873 36964 12877 37020
rect 12813 36960 12877 36964
rect 12893 37020 12957 37024
rect 12893 36964 12897 37020
rect 12897 36964 12953 37020
rect 12953 36964 12957 37020
rect 12893 36960 12957 36964
rect 12973 37020 13037 37024
rect 12973 36964 12977 37020
rect 12977 36964 13033 37020
rect 13033 36964 13037 37020
rect 12973 36960 13037 36964
rect 13053 37020 13117 37024
rect 13053 36964 13057 37020
rect 13057 36964 13113 37020
rect 13113 36964 13117 37020
rect 13053 36960 13117 36964
rect 3917 36476 3981 36480
rect 3917 36420 3921 36476
rect 3921 36420 3977 36476
rect 3977 36420 3981 36476
rect 3917 36416 3981 36420
rect 3997 36476 4061 36480
rect 3997 36420 4001 36476
rect 4001 36420 4057 36476
rect 4057 36420 4061 36476
rect 3997 36416 4061 36420
rect 4077 36476 4141 36480
rect 4077 36420 4081 36476
rect 4081 36420 4137 36476
rect 4137 36420 4141 36476
rect 4077 36416 4141 36420
rect 4157 36476 4221 36480
rect 4157 36420 4161 36476
rect 4161 36420 4217 36476
rect 4217 36420 4221 36476
rect 4157 36416 4221 36420
rect 9848 36476 9912 36480
rect 9848 36420 9852 36476
rect 9852 36420 9908 36476
rect 9908 36420 9912 36476
rect 9848 36416 9912 36420
rect 9928 36476 9992 36480
rect 9928 36420 9932 36476
rect 9932 36420 9988 36476
rect 9988 36420 9992 36476
rect 9928 36416 9992 36420
rect 10008 36476 10072 36480
rect 10008 36420 10012 36476
rect 10012 36420 10068 36476
rect 10068 36420 10072 36476
rect 10008 36416 10072 36420
rect 10088 36476 10152 36480
rect 10088 36420 10092 36476
rect 10092 36420 10148 36476
rect 10148 36420 10152 36476
rect 10088 36416 10152 36420
rect 15778 36476 15842 36480
rect 15778 36420 15782 36476
rect 15782 36420 15838 36476
rect 15838 36420 15842 36476
rect 15778 36416 15842 36420
rect 15858 36476 15922 36480
rect 15858 36420 15862 36476
rect 15862 36420 15918 36476
rect 15918 36420 15922 36476
rect 15858 36416 15922 36420
rect 15938 36476 16002 36480
rect 15938 36420 15942 36476
rect 15942 36420 15998 36476
rect 15998 36420 16002 36476
rect 15938 36416 16002 36420
rect 16018 36476 16082 36480
rect 16018 36420 16022 36476
rect 16022 36420 16078 36476
rect 16078 36420 16082 36476
rect 16018 36416 16082 36420
rect 6882 35932 6946 35936
rect 6882 35876 6886 35932
rect 6886 35876 6942 35932
rect 6942 35876 6946 35932
rect 6882 35872 6946 35876
rect 6962 35932 7026 35936
rect 6962 35876 6966 35932
rect 6966 35876 7022 35932
rect 7022 35876 7026 35932
rect 6962 35872 7026 35876
rect 7042 35932 7106 35936
rect 7042 35876 7046 35932
rect 7046 35876 7102 35932
rect 7102 35876 7106 35932
rect 7042 35872 7106 35876
rect 7122 35932 7186 35936
rect 7122 35876 7126 35932
rect 7126 35876 7182 35932
rect 7182 35876 7186 35932
rect 7122 35872 7186 35876
rect 12813 35932 12877 35936
rect 12813 35876 12817 35932
rect 12817 35876 12873 35932
rect 12873 35876 12877 35932
rect 12813 35872 12877 35876
rect 12893 35932 12957 35936
rect 12893 35876 12897 35932
rect 12897 35876 12953 35932
rect 12953 35876 12957 35932
rect 12893 35872 12957 35876
rect 12973 35932 13037 35936
rect 12973 35876 12977 35932
rect 12977 35876 13033 35932
rect 13033 35876 13037 35932
rect 12973 35872 13037 35876
rect 13053 35932 13117 35936
rect 13053 35876 13057 35932
rect 13057 35876 13113 35932
rect 13113 35876 13117 35932
rect 13053 35872 13117 35876
rect 3917 35388 3981 35392
rect 3917 35332 3921 35388
rect 3921 35332 3977 35388
rect 3977 35332 3981 35388
rect 3917 35328 3981 35332
rect 3997 35388 4061 35392
rect 3997 35332 4001 35388
rect 4001 35332 4057 35388
rect 4057 35332 4061 35388
rect 3997 35328 4061 35332
rect 4077 35388 4141 35392
rect 4077 35332 4081 35388
rect 4081 35332 4137 35388
rect 4137 35332 4141 35388
rect 4077 35328 4141 35332
rect 4157 35388 4221 35392
rect 4157 35332 4161 35388
rect 4161 35332 4217 35388
rect 4217 35332 4221 35388
rect 4157 35328 4221 35332
rect 9848 35388 9912 35392
rect 9848 35332 9852 35388
rect 9852 35332 9908 35388
rect 9908 35332 9912 35388
rect 9848 35328 9912 35332
rect 9928 35388 9992 35392
rect 9928 35332 9932 35388
rect 9932 35332 9988 35388
rect 9988 35332 9992 35388
rect 9928 35328 9992 35332
rect 10008 35388 10072 35392
rect 10008 35332 10012 35388
rect 10012 35332 10068 35388
rect 10068 35332 10072 35388
rect 10008 35328 10072 35332
rect 10088 35388 10152 35392
rect 10088 35332 10092 35388
rect 10092 35332 10148 35388
rect 10148 35332 10152 35388
rect 10088 35328 10152 35332
rect 15778 35388 15842 35392
rect 15778 35332 15782 35388
rect 15782 35332 15838 35388
rect 15838 35332 15842 35388
rect 15778 35328 15842 35332
rect 15858 35388 15922 35392
rect 15858 35332 15862 35388
rect 15862 35332 15918 35388
rect 15918 35332 15922 35388
rect 15858 35328 15922 35332
rect 15938 35388 16002 35392
rect 15938 35332 15942 35388
rect 15942 35332 15998 35388
rect 15998 35332 16002 35388
rect 15938 35328 16002 35332
rect 16018 35388 16082 35392
rect 16018 35332 16022 35388
rect 16022 35332 16078 35388
rect 16078 35332 16082 35388
rect 16018 35328 16082 35332
rect 6882 34844 6946 34848
rect 6882 34788 6886 34844
rect 6886 34788 6942 34844
rect 6942 34788 6946 34844
rect 6882 34784 6946 34788
rect 6962 34844 7026 34848
rect 6962 34788 6966 34844
rect 6966 34788 7022 34844
rect 7022 34788 7026 34844
rect 6962 34784 7026 34788
rect 7042 34844 7106 34848
rect 7042 34788 7046 34844
rect 7046 34788 7102 34844
rect 7102 34788 7106 34844
rect 7042 34784 7106 34788
rect 7122 34844 7186 34848
rect 7122 34788 7126 34844
rect 7126 34788 7182 34844
rect 7182 34788 7186 34844
rect 7122 34784 7186 34788
rect 12813 34844 12877 34848
rect 12813 34788 12817 34844
rect 12817 34788 12873 34844
rect 12873 34788 12877 34844
rect 12813 34784 12877 34788
rect 12893 34844 12957 34848
rect 12893 34788 12897 34844
rect 12897 34788 12953 34844
rect 12953 34788 12957 34844
rect 12893 34784 12957 34788
rect 12973 34844 13037 34848
rect 12973 34788 12977 34844
rect 12977 34788 13033 34844
rect 13033 34788 13037 34844
rect 12973 34784 13037 34788
rect 13053 34844 13117 34848
rect 13053 34788 13057 34844
rect 13057 34788 13113 34844
rect 13113 34788 13117 34844
rect 13053 34784 13117 34788
rect 3917 34300 3981 34304
rect 3917 34244 3921 34300
rect 3921 34244 3977 34300
rect 3977 34244 3981 34300
rect 3917 34240 3981 34244
rect 3997 34300 4061 34304
rect 3997 34244 4001 34300
rect 4001 34244 4057 34300
rect 4057 34244 4061 34300
rect 3997 34240 4061 34244
rect 4077 34300 4141 34304
rect 4077 34244 4081 34300
rect 4081 34244 4137 34300
rect 4137 34244 4141 34300
rect 4077 34240 4141 34244
rect 4157 34300 4221 34304
rect 4157 34244 4161 34300
rect 4161 34244 4217 34300
rect 4217 34244 4221 34300
rect 4157 34240 4221 34244
rect 9848 34300 9912 34304
rect 9848 34244 9852 34300
rect 9852 34244 9908 34300
rect 9908 34244 9912 34300
rect 9848 34240 9912 34244
rect 9928 34300 9992 34304
rect 9928 34244 9932 34300
rect 9932 34244 9988 34300
rect 9988 34244 9992 34300
rect 9928 34240 9992 34244
rect 10008 34300 10072 34304
rect 10008 34244 10012 34300
rect 10012 34244 10068 34300
rect 10068 34244 10072 34300
rect 10008 34240 10072 34244
rect 10088 34300 10152 34304
rect 10088 34244 10092 34300
rect 10092 34244 10148 34300
rect 10148 34244 10152 34300
rect 10088 34240 10152 34244
rect 15778 34300 15842 34304
rect 15778 34244 15782 34300
rect 15782 34244 15838 34300
rect 15838 34244 15842 34300
rect 15778 34240 15842 34244
rect 15858 34300 15922 34304
rect 15858 34244 15862 34300
rect 15862 34244 15918 34300
rect 15918 34244 15922 34300
rect 15858 34240 15922 34244
rect 15938 34300 16002 34304
rect 15938 34244 15942 34300
rect 15942 34244 15998 34300
rect 15998 34244 16002 34300
rect 15938 34240 16002 34244
rect 16018 34300 16082 34304
rect 16018 34244 16022 34300
rect 16022 34244 16078 34300
rect 16078 34244 16082 34300
rect 16018 34240 16082 34244
rect 6882 33756 6946 33760
rect 6882 33700 6886 33756
rect 6886 33700 6942 33756
rect 6942 33700 6946 33756
rect 6882 33696 6946 33700
rect 6962 33756 7026 33760
rect 6962 33700 6966 33756
rect 6966 33700 7022 33756
rect 7022 33700 7026 33756
rect 6962 33696 7026 33700
rect 7042 33756 7106 33760
rect 7042 33700 7046 33756
rect 7046 33700 7102 33756
rect 7102 33700 7106 33756
rect 7042 33696 7106 33700
rect 7122 33756 7186 33760
rect 7122 33700 7126 33756
rect 7126 33700 7182 33756
rect 7182 33700 7186 33756
rect 7122 33696 7186 33700
rect 12813 33756 12877 33760
rect 12813 33700 12817 33756
rect 12817 33700 12873 33756
rect 12873 33700 12877 33756
rect 12813 33696 12877 33700
rect 12893 33756 12957 33760
rect 12893 33700 12897 33756
rect 12897 33700 12953 33756
rect 12953 33700 12957 33756
rect 12893 33696 12957 33700
rect 12973 33756 13037 33760
rect 12973 33700 12977 33756
rect 12977 33700 13033 33756
rect 13033 33700 13037 33756
rect 12973 33696 13037 33700
rect 13053 33756 13117 33760
rect 13053 33700 13057 33756
rect 13057 33700 13113 33756
rect 13113 33700 13117 33756
rect 13053 33696 13117 33700
rect 3917 33212 3981 33216
rect 3917 33156 3921 33212
rect 3921 33156 3977 33212
rect 3977 33156 3981 33212
rect 3917 33152 3981 33156
rect 3997 33212 4061 33216
rect 3997 33156 4001 33212
rect 4001 33156 4057 33212
rect 4057 33156 4061 33212
rect 3997 33152 4061 33156
rect 4077 33212 4141 33216
rect 4077 33156 4081 33212
rect 4081 33156 4137 33212
rect 4137 33156 4141 33212
rect 4077 33152 4141 33156
rect 4157 33212 4221 33216
rect 4157 33156 4161 33212
rect 4161 33156 4217 33212
rect 4217 33156 4221 33212
rect 4157 33152 4221 33156
rect 9848 33212 9912 33216
rect 9848 33156 9852 33212
rect 9852 33156 9908 33212
rect 9908 33156 9912 33212
rect 9848 33152 9912 33156
rect 9928 33212 9992 33216
rect 9928 33156 9932 33212
rect 9932 33156 9988 33212
rect 9988 33156 9992 33212
rect 9928 33152 9992 33156
rect 10008 33212 10072 33216
rect 10008 33156 10012 33212
rect 10012 33156 10068 33212
rect 10068 33156 10072 33212
rect 10008 33152 10072 33156
rect 10088 33212 10152 33216
rect 10088 33156 10092 33212
rect 10092 33156 10148 33212
rect 10148 33156 10152 33212
rect 10088 33152 10152 33156
rect 15778 33212 15842 33216
rect 15778 33156 15782 33212
rect 15782 33156 15838 33212
rect 15838 33156 15842 33212
rect 15778 33152 15842 33156
rect 15858 33212 15922 33216
rect 15858 33156 15862 33212
rect 15862 33156 15918 33212
rect 15918 33156 15922 33212
rect 15858 33152 15922 33156
rect 15938 33212 16002 33216
rect 15938 33156 15942 33212
rect 15942 33156 15998 33212
rect 15998 33156 16002 33212
rect 15938 33152 16002 33156
rect 16018 33212 16082 33216
rect 16018 33156 16022 33212
rect 16022 33156 16078 33212
rect 16078 33156 16082 33212
rect 16018 33152 16082 33156
rect 6882 32668 6946 32672
rect 6882 32612 6886 32668
rect 6886 32612 6942 32668
rect 6942 32612 6946 32668
rect 6882 32608 6946 32612
rect 6962 32668 7026 32672
rect 6962 32612 6966 32668
rect 6966 32612 7022 32668
rect 7022 32612 7026 32668
rect 6962 32608 7026 32612
rect 7042 32668 7106 32672
rect 7042 32612 7046 32668
rect 7046 32612 7102 32668
rect 7102 32612 7106 32668
rect 7042 32608 7106 32612
rect 7122 32668 7186 32672
rect 7122 32612 7126 32668
rect 7126 32612 7182 32668
rect 7182 32612 7186 32668
rect 7122 32608 7186 32612
rect 12813 32668 12877 32672
rect 12813 32612 12817 32668
rect 12817 32612 12873 32668
rect 12873 32612 12877 32668
rect 12813 32608 12877 32612
rect 12893 32668 12957 32672
rect 12893 32612 12897 32668
rect 12897 32612 12953 32668
rect 12953 32612 12957 32668
rect 12893 32608 12957 32612
rect 12973 32668 13037 32672
rect 12973 32612 12977 32668
rect 12977 32612 13033 32668
rect 13033 32612 13037 32668
rect 12973 32608 13037 32612
rect 13053 32668 13117 32672
rect 13053 32612 13057 32668
rect 13057 32612 13113 32668
rect 13113 32612 13117 32668
rect 13053 32608 13117 32612
rect 3917 32124 3981 32128
rect 3917 32068 3921 32124
rect 3921 32068 3977 32124
rect 3977 32068 3981 32124
rect 3917 32064 3981 32068
rect 3997 32124 4061 32128
rect 3997 32068 4001 32124
rect 4001 32068 4057 32124
rect 4057 32068 4061 32124
rect 3997 32064 4061 32068
rect 4077 32124 4141 32128
rect 4077 32068 4081 32124
rect 4081 32068 4137 32124
rect 4137 32068 4141 32124
rect 4077 32064 4141 32068
rect 4157 32124 4221 32128
rect 4157 32068 4161 32124
rect 4161 32068 4217 32124
rect 4217 32068 4221 32124
rect 4157 32064 4221 32068
rect 9848 32124 9912 32128
rect 9848 32068 9852 32124
rect 9852 32068 9908 32124
rect 9908 32068 9912 32124
rect 9848 32064 9912 32068
rect 9928 32124 9992 32128
rect 9928 32068 9932 32124
rect 9932 32068 9988 32124
rect 9988 32068 9992 32124
rect 9928 32064 9992 32068
rect 10008 32124 10072 32128
rect 10008 32068 10012 32124
rect 10012 32068 10068 32124
rect 10068 32068 10072 32124
rect 10008 32064 10072 32068
rect 10088 32124 10152 32128
rect 10088 32068 10092 32124
rect 10092 32068 10148 32124
rect 10148 32068 10152 32124
rect 10088 32064 10152 32068
rect 15778 32124 15842 32128
rect 15778 32068 15782 32124
rect 15782 32068 15838 32124
rect 15838 32068 15842 32124
rect 15778 32064 15842 32068
rect 15858 32124 15922 32128
rect 15858 32068 15862 32124
rect 15862 32068 15918 32124
rect 15918 32068 15922 32124
rect 15858 32064 15922 32068
rect 15938 32124 16002 32128
rect 15938 32068 15942 32124
rect 15942 32068 15998 32124
rect 15998 32068 16002 32124
rect 15938 32064 16002 32068
rect 16018 32124 16082 32128
rect 16018 32068 16022 32124
rect 16022 32068 16078 32124
rect 16078 32068 16082 32124
rect 16018 32064 16082 32068
rect 6882 31580 6946 31584
rect 6882 31524 6886 31580
rect 6886 31524 6942 31580
rect 6942 31524 6946 31580
rect 6882 31520 6946 31524
rect 6962 31580 7026 31584
rect 6962 31524 6966 31580
rect 6966 31524 7022 31580
rect 7022 31524 7026 31580
rect 6962 31520 7026 31524
rect 7042 31580 7106 31584
rect 7042 31524 7046 31580
rect 7046 31524 7102 31580
rect 7102 31524 7106 31580
rect 7042 31520 7106 31524
rect 7122 31580 7186 31584
rect 7122 31524 7126 31580
rect 7126 31524 7182 31580
rect 7182 31524 7186 31580
rect 7122 31520 7186 31524
rect 12813 31580 12877 31584
rect 12813 31524 12817 31580
rect 12817 31524 12873 31580
rect 12873 31524 12877 31580
rect 12813 31520 12877 31524
rect 12893 31580 12957 31584
rect 12893 31524 12897 31580
rect 12897 31524 12953 31580
rect 12953 31524 12957 31580
rect 12893 31520 12957 31524
rect 12973 31580 13037 31584
rect 12973 31524 12977 31580
rect 12977 31524 13033 31580
rect 13033 31524 13037 31580
rect 12973 31520 13037 31524
rect 13053 31580 13117 31584
rect 13053 31524 13057 31580
rect 13057 31524 13113 31580
rect 13113 31524 13117 31580
rect 13053 31520 13117 31524
rect 3917 31036 3981 31040
rect 3917 30980 3921 31036
rect 3921 30980 3977 31036
rect 3977 30980 3981 31036
rect 3917 30976 3981 30980
rect 3997 31036 4061 31040
rect 3997 30980 4001 31036
rect 4001 30980 4057 31036
rect 4057 30980 4061 31036
rect 3997 30976 4061 30980
rect 4077 31036 4141 31040
rect 4077 30980 4081 31036
rect 4081 30980 4137 31036
rect 4137 30980 4141 31036
rect 4077 30976 4141 30980
rect 4157 31036 4221 31040
rect 4157 30980 4161 31036
rect 4161 30980 4217 31036
rect 4217 30980 4221 31036
rect 4157 30976 4221 30980
rect 9848 31036 9912 31040
rect 9848 30980 9852 31036
rect 9852 30980 9908 31036
rect 9908 30980 9912 31036
rect 9848 30976 9912 30980
rect 9928 31036 9992 31040
rect 9928 30980 9932 31036
rect 9932 30980 9988 31036
rect 9988 30980 9992 31036
rect 9928 30976 9992 30980
rect 10008 31036 10072 31040
rect 10008 30980 10012 31036
rect 10012 30980 10068 31036
rect 10068 30980 10072 31036
rect 10008 30976 10072 30980
rect 10088 31036 10152 31040
rect 10088 30980 10092 31036
rect 10092 30980 10148 31036
rect 10148 30980 10152 31036
rect 10088 30976 10152 30980
rect 15778 31036 15842 31040
rect 15778 30980 15782 31036
rect 15782 30980 15838 31036
rect 15838 30980 15842 31036
rect 15778 30976 15842 30980
rect 15858 31036 15922 31040
rect 15858 30980 15862 31036
rect 15862 30980 15918 31036
rect 15918 30980 15922 31036
rect 15858 30976 15922 30980
rect 15938 31036 16002 31040
rect 15938 30980 15942 31036
rect 15942 30980 15998 31036
rect 15998 30980 16002 31036
rect 15938 30976 16002 30980
rect 16018 31036 16082 31040
rect 16018 30980 16022 31036
rect 16022 30980 16078 31036
rect 16078 30980 16082 31036
rect 16018 30976 16082 30980
rect 6882 30492 6946 30496
rect 6882 30436 6886 30492
rect 6886 30436 6942 30492
rect 6942 30436 6946 30492
rect 6882 30432 6946 30436
rect 6962 30492 7026 30496
rect 6962 30436 6966 30492
rect 6966 30436 7022 30492
rect 7022 30436 7026 30492
rect 6962 30432 7026 30436
rect 7042 30492 7106 30496
rect 7042 30436 7046 30492
rect 7046 30436 7102 30492
rect 7102 30436 7106 30492
rect 7042 30432 7106 30436
rect 7122 30492 7186 30496
rect 7122 30436 7126 30492
rect 7126 30436 7182 30492
rect 7182 30436 7186 30492
rect 7122 30432 7186 30436
rect 12813 30492 12877 30496
rect 12813 30436 12817 30492
rect 12817 30436 12873 30492
rect 12873 30436 12877 30492
rect 12813 30432 12877 30436
rect 12893 30492 12957 30496
rect 12893 30436 12897 30492
rect 12897 30436 12953 30492
rect 12953 30436 12957 30492
rect 12893 30432 12957 30436
rect 12973 30492 13037 30496
rect 12973 30436 12977 30492
rect 12977 30436 13033 30492
rect 13033 30436 13037 30492
rect 12973 30432 13037 30436
rect 13053 30492 13117 30496
rect 13053 30436 13057 30492
rect 13057 30436 13113 30492
rect 13113 30436 13117 30492
rect 13053 30432 13117 30436
rect 3917 29948 3981 29952
rect 3917 29892 3921 29948
rect 3921 29892 3977 29948
rect 3977 29892 3981 29948
rect 3917 29888 3981 29892
rect 3997 29948 4061 29952
rect 3997 29892 4001 29948
rect 4001 29892 4057 29948
rect 4057 29892 4061 29948
rect 3997 29888 4061 29892
rect 4077 29948 4141 29952
rect 4077 29892 4081 29948
rect 4081 29892 4137 29948
rect 4137 29892 4141 29948
rect 4077 29888 4141 29892
rect 4157 29948 4221 29952
rect 4157 29892 4161 29948
rect 4161 29892 4217 29948
rect 4217 29892 4221 29948
rect 4157 29888 4221 29892
rect 9848 29948 9912 29952
rect 9848 29892 9852 29948
rect 9852 29892 9908 29948
rect 9908 29892 9912 29948
rect 9848 29888 9912 29892
rect 9928 29948 9992 29952
rect 9928 29892 9932 29948
rect 9932 29892 9988 29948
rect 9988 29892 9992 29948
rect 9928 29888 9992 29892
rect 10008 29948 10072 29952
rect 10008 29892 10012 29948
rect 10012 29892 10068 29948
rect 10068 29892 10072 29948
rect 10008 29888 10072 29892
rect 10088 29948 10152 29952
rect 10088 29892 10092 29948
rect 10092 29892 10148 29948
rect 10148 29892 10152 29948
rect 10088 29888 10152 29892
rect 15778 29948 15842 29952
rect 15778 29892 15782 29948
rect 15782 29892 15838 29948
rect 15838 29892 15842 29948
rect 15778 29888 15842 29892
rect 15858 29948 15922 29952
rect 15858 29892 15862 29948
rect 15862 29892 15918 29948
rect 15918 29892 15922 29948
rect 15858 29888 15922 29892
rect 15938 29948 16002 29952
rect 15938 29892 15942 29948
rect 15942 29892 15998 29948
rect 15998 29892 16002 29948
rect 15938 29888 16002 29892
rect 16018 29948 16082 29952
rect 16018 29892 16022 29948
rect 16022 29892 16078 29948
rect 16078 29892 16082 29948
rect 16018 29888 16082 29892
rect 6882 29404 6946 29408
rect 6882 29348 6886 29404
rect 6886 29348 6942 29404
rect 6942 29348 6946 29404
rect 6882 29344 6946 29348
rect 6962 29404 7026 29408
rect 6962 29348 6966 29404
rect 6966 29348 7022 29404
rect 7022 29348 7026 29404
rect 6962 29344 7026 29348
rect 7042 29404 7106 29408
rect 7042 29348 7046 29404
rect 7046 29348 7102 29404
rect 7102 29348 7106 29404
rect 7042 29344 7106 29348
rect 7122 29404 7186 29408
rect 7122 29348 7126 29404
rect 7126 29348 7182 29404
rect 7182 29348 7186 29404
rect 7122 29344 7186 29348
rect 12813 29404 12877 29408
rect 12813 29348 12817 29404
rect 12817 29348 12873 29404
rect 12873 29348 12877 29404
rect 12813 29344 12877 29348
rect 12893 29404 12957 29408
rect 12893 29348 12897 29404
rect 12897 29348 12953 29404
rect 12953 29348 12957 29404
rect 12893 29344 12957 29348
rect 12973 29404 13037 29408
rect 12973 29348 12977 29404
rect 12977 29348 13033 29404
rect 13033 29348 13037 29404
rect 12973 29344 13037 29348
rect 13053 29404 13117 29408
rect 13053 29348 13057 29404
rect 13057 29348 13113 29404
rect 13113 29348 13117 29404
rect 13053 29344 13117 29348
rect 3917 28860 3981 28864
rect 3917 28804 3921 28860
rect 3921 28804 3977 28860
rect 3977 28804 3981 28860
rect 3917 28800 3981 28804
rect 3997 28860 4061 28864
rect 3997 28804 4001 28860
rect 4001 28804 4057 28860
rect 4057 28804 4061 28860
rect 3997 28800 4061 28804
rect 4077 28860 4141 28864
rect 4077 28804 4081 28860
rect 4081 28804 4137 28860
rect 4137 28804 4141 28860
rect 4077 28800 4141 28804
rect 4157 28860 4221 28864
rect 4157 28804 4161 28860
rect 4161 28804 4217 28860
rect 4217 28804 4221 28860
rect 4157 28800 4221 28804
rect 9848 28860 9912 28864
rect 9848 28804 9852 28860
rect 9852 28804 9908 28860
rect 9908 28804 9912 28860
rect 9848 28800 9912 28804
rect 9928 28860 9992 28864
rect 9928 28804 9932 28860
rect 9932 28804 9988 28860
rect 9988 28804 9992 28860
rect 9928 28800 9992 28804
rect 10008 28860 10072 28864
rect 10008 28804 10012 28860
rect 10012 28804 10068 28860
rect 10068 28804 10072 28860
rect 10008 28800 10072 28804
rect 10088 28860 10152 28864
rect 10088 28804 10092 28860
rect 10092 28804 10148 28860
rect 10148 28804 10152 28860
rect 10088 28800 10152 28804
rect 15778 28860 15842 28864
rect 15778 28804 15782 28860
rect 15782 28804 15838 28860
rect 15838 28804 15842 28860
rect 15778 28800 15842 28804
rect 15858 28860 15922 28864
rect 15858 28804 15862 28860
rect 15862 28804 15918 28860
rect 15918 28804 15922 28860
rect 15858 28800 15922 28804
rect 15938 28860 16002 28864
rect 15938 28804 15942 28860
rect 15942 28804 15998 28860
rect 15998 28804 16002 28860
rect 15938 28800 16002 28804
rect 16018 28860 16082 28864
rect 16018 28804 16022 28860
rect 16022 28804 16078 28860
rect 16078 28804 16082 28860
rect 16018 28800 16082 28804
rect 6882 28316 6946 28320
rect 6882 28260 6886 28316
rect 6886 28260 6942 28316
rect 6942 28260 6946 28316
rect 6882 28256 6946 28260
rect 6962 28316 7026 28320
rect 6962 28260 6966 28316
rect 6966 28260 7022 28316
rect 7022 28260 7026 28316
rect 6962 28256 7026 28260
rect 7042 28316 7106 28320
rect 7042 28260 7046 28316
rect 7046 28260 7102 28316
rect 7102 28260 7106 28316
rect 7042 28256 7106 28260
rect 7122 28316 7186 28320
rect 7122 28260 7126 28316
rect 7126 28260 7182 28316
rect 7182 28260 7186 28316
rect 7122 28256 7186 28260
rect 12813 28316 12877 28320
rect 12813 28260 12817 28316
rect 12817 28260 12873 28316
rect 12873 28260 12877 28316
rect 12813 28256 12877 28260
rect 12893 28316 12957 28320
rect 12893 28260 12897 28316
rect 12897 28260 12953 28316
rect 12953 28260 12957 28316
rect 12893 28256 12957 28260
rect 12973 28316 13037 28320
rect 12973 28260 12977 28316
rect 12977 28260 13033 28316
rect 13033 28260 13037 28316
rect 12973 28256 13037 28260
rect 13053 28316 13117 28320
rect 13053 28260 13057 28316
rect 13057 28260 13113 28316
rect 13113 28260 13117 28316
rect 13053 28256 13117 28260
rect 3917 27772 3981 27776
rect 3917 27716 3921 27772
rect 3921 27716 3977 27772
rect 3977 27716 3981 27772
rect 3917 27712 3981 27716
rect 3997 27772 4061 27776
rect 3997 27716 4001 27772
rect 4001 27716 4057 27772
rect 4057 27716 4061 27772
rect 3997 27712 4061 27716
rect 4077 27772 4141 27776
rect 4077 27716 4081 27772
rect 4081 27716 4137 27772
rect 4137 27716 4141 27772
rect 4077 27712 4141 27716
rect 4157 27772 4221 27776
rect 4157 27716 4161 27772
rect 4161 27716 4217 27772
rect 4217 27716 4221 27772
rect 4157 27712 4221 27716
rect 9848 27772 9912 27776
rect 9848 27716 9852 27772
rect 9852 27716 9908 27772
rect 9908 27716 9912 27772
rect 9848 27712 9912 27716
rect 9928 27772 9992 27776
rect 9928 27716 9932 27772
rect 9932 27716 9988 27772
rect 9988 27716 9992 27772
rect 9928 27712 9992 27716
rect 10008 27772 10072 27776
rect 10008 27716 10012 27772
rect 10012 27716 10068 27772
rect 10068 27716 10072 27772
rect 10008 27712 10072 27716
rect 10088 27772 10152 27776
rect 10088 27716 10092 27772
rect 10092 27716 10148 27772
rect 10148 27716 10152 27772
rect 10088 27712 10152 27716
rect 15778 27772 15842 27776
rect 15778 27716 15782 27772
rect 15782 27716 15838 27772
rect 15838 27716 15842 27772
rect 15778 27712 15842 27716
rect 15858 27772 15922 27776
rect 15858 27716 15862 27772
rect 15862 27716 15918 27772
rect 15918 27716 15922 27772
rect 15858 27712 15922 27716
rect 15938 27772 16002 27776
rect 15938 27716 15942 27772
rect 15942 27716 15998 27772
rect 15998 27716 16002 27772
rect 15938 27712 16002 27716
rect 16018 27772 16082 27776
rect 16018 27716 16022 27772
rect 16022 27716 16078 27772
rect 16078 27716 16082 27772
rect 16018 27712 16082 27716
rect 6882 27228 6946 27232
rect 6882 27172 6886 27228
rect 6886 27172 6942 27228
rect 6942 27172 6946 27228
rect 6882 27168 6946 27172
rect 6962 27228 7026 27232
rect 6962 27172 6966 27228
rect 6966 27172 7022 27228
rect 7022 27172 7026 27228
rect 6962 27168 7026 27172
rect 7042 27228 7106 27232
rect 7042 27172 7046 27228
rect 7046 27172 7102 27228
rect 7102 27172 7106 27228
rect 7042 27168 7106 27172
rect 7122 27228 7186 27232
rect 7122 27172 7126 27228
rect 7126 27172 7182 27228
rect 7182 27172 7186 27228
rect 7122 27168 7186 27172
rect 12813 27228 12877 27232
rect 12813 27172 12817 27228
rect 12817 27172 12873 27228
rect 12873 27172 12877 27228
rect 12813 27168 12877 27172
rect 12893 27228 12957 27232
rect 12893 27172 12897 27228
rect 12897 27172 12953 27228
rect 12953 27172 12957 27228
rect 12893 27168 12957 27172
rect 12973 27228 13037 27232
rect 12973 27172 12977 27228
rect 12977 27172 13033 27228
rect 13033 27172 13037 27228
rect 12973 27168 13037 27172
rect 13053 27228 13117 27232
rect 13053 27172 13057 27228
rect 13057 27172 13113 27228
rect 13113 27172 13117 27228
rect 13053 27168 13117 27172
rect 3917 26684 3981 26688
rect 3917 26628 3921 26684
rect 3921 26628 3977 26684
rect 3977 26628 3981 26684
rect 3917 26624 3981 26628
rect 3997 26684 4061 26688
rect 3997 26628 4001 26684
rect 4001 26628 4057 26684
rect 4057 26628 4061 26684
rect 3997 26624 4061 26628
rect 4077 26684 4141 26688
rect 4077 26628 4081 26684
rect 4081 26628 4137 26684
rect 4137 26628 4141 26684
rect 4077 26624 4141 26628
rect 4157 26684 4221 26688
rect 4157 26628 4161 26684
rect 4161 26628 4217 26684
rect 4217 26628 4221 26684
rect 4157 26624 4221 26628
rect 9848 26684 9912 26688
rect 9848 26628 9852 26684
rect 9852 26628 9908 26684
rect 9908 26628 9912 26684
rect 9848 26624 9912 26628
rect 9928 26684 9992 26688
rect 9928 26628 9932 26684
rect 9932 26628 9988 26684
rect 9988 26628 9992 26684
rect 9928 26624 9992 26628
rect 10008 26684 10072 26688
rect 10008 26628 10012 26684
rect 10012 26628 10068 26684
rect 10068 26628 10072 26684
rect 10008 26624 10072 26628
rect 10088 26684 10152 26688
rect 10088 26628 10092 26684
rect 10092 26628 10148 26684
rect 10148 26628 10152 26684
rect 10088 26624 10152 26628
rect 15778 26684 15842 26688
rect 15778 26628 15782 26684
rect 15782 26628 15838 26684
rect 15838 26628 15842 26684
rect 15778 26624 15842 26628
rect 15858 26684 15922 26688
rect 15858 26628 15862 26684
rect 15862 26628 15918 26684
rect 15918 26628 15922 26684
rect 15858 26624 15922 26628
rect 15938 26684 16002 26688
rect 15938 26628 15942 26684
rect 15942 26628 15998 26684
rect 15998 26628 16002 26684
rect 15938 26624 16002 26628
rect 16018 26684 16082 26688
rect 16018 26628 16022 26684
rect 16022 26628 16078 26684
rect 16078 26628 16082 26684
rect 16018 26624 16082 26628
rect 6882 26140 6946 26144
rect 6882 26084 6886 26140
rect 6886 26084 6942 26140
rect 6942 26084 6946 26140
rect 6882 26080 6946 26084
rect 6962 26140 7026 26144
rect 6962 26084 6966 26140
rect 6966 26084 7022 26140
rect 7022 26084 7026 26140
rect 6962 26080 7026 26084
rect 7042 26140 7106 26144
rect 7042 26084 7046 26140
rect 7046 26084 7102 26140
rect 7102 26084 7106 26140
rect 7042 26080 7106 26084
rect 7122 26140 7186 26144
rect 7122 26084 7126 26140
rect 7126 26084 7182 26140
rect 7182 26084 7186 26140
rect 7122 26080 7186 26084
rect 12813 26140 12877 26144
rect 12813 26084 12817 26140
rect 12817 26084 12873 26140
rect 12873 26084 12877 26140
rect 12813 26080 12877 26084
rect 12893 26140 12957 26144
rect 12893 26084 12897 26140
rect 12897 26084 12953 26140
rect 12953 26084 12957 26140
rect 12893 26080 12957 26084
rect 12973 26140 13037 26144
rect 12973 26084 12977 26140
rect 12977 26084 13033 26140
rect 13033 26084 13037 26140
rect 12973 26080 13037 26084
rect 13053 26140 13117 26144
rect 13053 26084 13057 26140
rect 13057 26084 13113 26140
rect 13113 26084 13117 26140
rect 13053 26080 13117 26084
rect 3917 25596 3981 25600
rect 3917 25540 3921 25596
rect 3921 25540 3977 25596
rect 3977 25540 3981 25596
rect 3917 25536 3981 25540
rect 3997 25596 4061 25600
rect 3997 25540 4001 25596
rect 4001 25540 4057 25596
rect 4057 25540 4061 25596
rect 3997 25536 4061 25540
rect 4077 25596 4141 25600
rect 4077 25540 4081 25596
rect 4081 25540 4137 25596
rect 4137 25540 4141 25596
rect 4077 25536 4141 25540
rect 4157 25596 4221 25600
rect 4157 25540 4161 25596
rect 4161 25540 4217 25596
rect 4217 25540 4221 25596
rect 4157 25536 4221 25540
rect 9848 25596 9912 25600
rect 9848 25540 9852 25596
rect 9852 25540 9908 25596
rect 9908 25540 9912 25596
rect 9848 25536 9912 25540
rect 9928 25596 9992 25600
rect 9928 25540 9932 25596
rect 9932 25540 9988 25596
rect 9988 25540 9992 25596
rect 9928 25536 9992 25540
rect 10008 25596 10072 25600
rect 10008 25540 10012 25596
rect 10012 25540 10068 25596
rect 10068 25540 10072 25596
rect 10008 25536 10072 25540
rect 10088 25596 10152 25600
rect 10088 25540 10092 25596
rect 10092 25540 10148 25596
rect 10148 25540 10152 25596
rect 10088 25536 10152 25540
rect 15778 25596 15842 25600
rect 15778 25540 15782 25596
rect 15782 25540 15838 25596
rect 15838 25540 15842 25596
rect 15778 25536 15842 25540
rect 15858 25596 15922 25600
rect 15858 25540 15862 25596
rect 15862 25540 15918 25596
rect 15918 25540 15922 25596
rect 15858 25536 15922 25540
rect 15938 25596 16002 25600
rect 15938 25540 15942 25596
rect 15942 25540 15998 25596
rect 15998 25540 16002 25596
rect 15938 25536 16002 25540
rect 16018 25596 16082 25600
rect 16018 25540 16022 25596
rect 16022 25540 16078 25596
rect 16078 25540 16082 25596
rect 16018 25536 16082 25540
rect 6882 25052 6946 25056
rect 6882 24996 6886 25052
rect 6886 24996 6942 25052
rect 6942 24996 6946 25052
rect 6882 24992 6946 24996
rect 6962 25052 7026 25056
rect 6962 24996 6966 25052
rect 6966 24996 7022 25052
rect 7022 24996 7026 25052
rect 6962 24992 7026 24996
rect 7042 25052 7106 25056
rect 7042 24996 7046 25052
rect 7046 24996 7102 25052
rect 7102 24996 7106 25052
rect 7042 24992 7106 24996
rect 7122 25052 7186 25056
rect 7122 24996 7126 25052
rect 7126 24996 7182 25052
rect 7182 24996 7186 25052
rect 7122 24992 7186 24996
rect 12813 25052 12877 25056
rect 12813 24996 12817 25052
rect 12817 24996 12873 25052
rect 12873 24996 12877 25052
rect 12813 24992 12877 24996
rect 12893 25052 12957 25056
rect 12893 24996 12897 25052
rect 12897 24996 12953 25052
rect 12953 24996 12957 25052
rect 12893 24992 12957 24996
rect 12973 25052 13037 25056
rect 12973 24996 12977 25052
rect 12977 24996 13033 25052
rect 13033 24996 13037 25052
rect 12973 24992 13037 24996
rect 13053 25052 13117 25056
rect 13053 24996 13057 25052
rect 13057 24996 13113 25052
rect 13113 24996 13117 25052
rect 13053 24992 13117 24996
rect 3917 24508 3981 24512
rect 3917 24452 3921 24508
rect 3921 24452 3977 24508
rect 3977 24452 3981 24508
rect 3917 24448 3981 24452
rect 3997 24508 4061 24512
rect 3997 24452 4001 24508
rect 4001 24452 4057 24508
rect 4057 24452 4061 24508
rect 3997 24448 4061 24452
rect 4077 24508 4141 24512
rect 4077 24452 4081 24508
rect 4081 24452 4137 24508
rect 4137 24452 4141 24508
rect 4077 24448 4141 24452
rect 4157 24508 4221 24512
rect 4157 24452 4161 24508
rect 4161 24452 4217 24508
rect 4217 24452 4221 24508
rect 4157 24448 4221 24452
rect 9848 24508 9912 24512
rect 9848 24452 9852 24508
rect 9852 24452 9908 24508
rect 9908 24452 9912 24508
rect 9848 24448 9912 24452
rect 9928 24508 9992 24512
rect 9928 24452 9932 24508
rect 9932 24452 9988 24508
rect 9988 24452 9992 24508
rect 9928 24448 9992 24452
rect 10008 24508 10072 24512
rect 10008 24452 10012 24508
rect 10012 24452 10068 24508
rect 10068 24452 10072 24508
rect 10008 24448 10072 24452
rect 10088 24508 10152 24512
rect 10088 24452 10092 24508
rect 10092 24452 10148 24508
rect 10148 24452 10152 24508
rect 10088 24448 10152 24452
rect 15778 24508 15842 24512
rect 15778 24452 15782 24508
rect 15782 24452 15838 24508
rect 15838 24452 15842 24508
rect 15778 24448 15842 24452
rect 15858 24508 15922 24512
rect 15858 24452 15862 24508
rect 15862 24452 15918 24508
rect 15918 24452 15922 24508
rect 15858 24448 15922 24452
rect 15938 24508 16002 24512
rect 15938 24452 15942 24508
rect 15942 24452 15998 24508
rect 15998 24452 16002 24508
rect 15938 24448 16002 24452
rect 16018 24508 16082 24512
rect 16018 24452 16022 24508
rect 16022 24452 16078 24508
rect 16078 24452 16082 24508
rect 16018 24448 16082 24452
rect 6882 23964 6946 23968
rect 6882 23908 6886 23964
rect 6886 23908 6942 23964
rect 6942 23908 6946 23964
rect 6882 23904 6946 23908
rect 6962 23964 7026 23968
rect 6962 23908 6966 23964
rect 6966 23908 7022 23964
rect 7022 23908 7026 23964
rect 6962 23904 7026 23908
rect 7042 23964 7106 23968
rect 7042 23908 7046 23964
rect 7046 23908 7102 23964
rect 7102 23908 7106 23964
rect 7042 23904 7106 23908
rect 7122 23964 7186 23968
rect 7122 23908 7126 23964
rect 7126 23908 7182 23964
rect 7182 23908 7186 23964
rect 7122 23904 7186 23908
rect 12813 23964 12877 23968
rect 12813 23908 12817 23964
rect 12817 23908 12873 23964
rect 12873 23908 12877 23964
rect 12813 23904 12877 23908
rect 12893 23964 12957 23968
rect 12893 23908 12897 23964
rect 12897 23908 12953 23964
rect 12953 23908 12957 23964
rect 12893 23904 12957 23908
rect 12973 23964 13037 23968
rect 12973 23908 12977 23964
rect 12977 23908 13033 23964
rect 13033 23908 13037 23964
rect 12973 23904 13037 23908
rect 13053 23964 13117 23968
rect 13053 23908 13057 23964
rect 13057 23908 13113 23964
rect 13113 23908 13117 23964
rect 13053 23904 13117 23908
rect 3917 23420 3981 23424
rect 3917 23364 3921 23420
rect 3921 23364 3977 23420
rect 3977 23364 3981 23420
rect 3917 23360 3981 23364
rect 3997 23420 4061 23424
rect 3997 23364 4001 23420
rect 4001 23364 4057 23420
rect 4057 23364 4061 23420
rect 3997 23360 4061 23364
rect 4077 23420 4141 23424
rect 4077 23364 4081 23420
rect 4081 23364 4137 23420
rect 4137 23364 4141 23420
rect 4077 23360 4141 23364
rect 4157 23420 4221 23424
rect 4157 23364 4161 23420
rect 4161 23364 4217 23420
rect 4217 23364 4221 23420
rect 4157 23360 4221 23364
rect 9848 23420 9912 23424
rect 9848 23364 9852 23420
rect 9852 23364 9908 23420
rect 9908 23364 9912 23420
rect 9848 23360 9912 23364
rect 9928 23420 9992 23424
rect 9928 23364 9932 23420
rect 9932 23364 9988 23420
rect 9988 23364 9992 23420
rect 9928 23360 9992 23364
rect 10008 23420 10072 23424
rect 10008 23364 10012 23420
rect 10012 23364 10068 23420
rect 10068 23364 10072 23420
rect 10008 23360 10072 23364
rect 10088 23420 10152 23424
rect 10088 23364 10092 23420
rect 10092 23364 10148 23420
rect 10148 23364 10152 23420
rect 10088 23360 10152 23364
rect 15778 23420 15842 23424
rect 15778 23364 15782 23420
rect 15782 23364 15838 23420
rect 15838 23364 15842 23420
rect 15778 23360 15842 23364
rect 15858 23420 15922 23424
rect 15858 23364 15862 23420
rect 15862 23364 15918 23420
rect 15918 23364 15922 23420
rect 15858 23360 15922 23364
rect 15938 23420 16002 23424
rect 15938 23364 15942 23420
rect 15942 23364 15998 23420
rect 15998 23364 16002 23420
rect 15938 23360 16002 23364
rect 16018 23420 16082 23424
rect 16018 23364 16022 23420
rect 16022 23364 16078 23420
rect 16078 23364 16082 23420
rect 16018 23360 16082 23364
rect 6882 22876 6946 22880
rect 6882 22820 6886 22876
rect 6886 22820 6942 22876
rect 6942 22820 6946 22876
rect 6882 22816 6946 22820
rect 6962 22876 7026 22880
rect 6962 22820 6966 22876
rect 6966 22820 7022 22876
rect 7022 22820 7026 22876
rect 6962 22816 7026 22820
rect 7042 22876 7106 22880
rect 7042 22820 7046 22876
rect 7046 22820 7102 22876
rect 7102 22820 7106 22876
rect 7042 22816 7106 22820
rect 7122 22876 7186 22880
rect 7122 22820 7126 22876
rect 7126 22820 7182 22876
rect 7182 22820 7186 22876
rect 7122 22816 7186 22820
rect 12813 22876 12877 22880
rect 12813 22820 12817 22876
rect 12817 22820 12873 22876
rect 12873 22820 12877 22876
rect 12813 22816 12877 22820
rect 12893 22876 12957 22880
rect 12893 22820 12897 22876
rect 12897 22820 12953 22876
rect 12953 22820 12957 22876
rect 12893 22816 12957 22820
rect 12973 22876 13037 22880
rect 12973 22820 12977 22876
rect 12977 22820 13033 22876
rect 13033 22820 13037 22876
rect 12973 22816 13037 22820
rect 13053 22876 13117 22880
rect 13053 22820 13057 22876
rect 13057 22820 13113 22876
rect 13113 22820 13117 22876
rect 13053 22816 13117 22820
rect 3917 22332 3981 22336
rect 3917 22276 3921 22332
rect 3921 22276 3977 22332
rect 3977 22276 3981 22332
rect 3917 22272 3981 22276
rect 3997 22332 4061 22336
rect 3997 22276 4001 22332
rect 4001 22276 4057 22332
rect 4057 22276 4061 22332
rect 3997 22272 4061 22276
rect 4077 22332 4141 22336
rect 4077 22276 4081 22332
rect 4081 22276 4137 22332
rect 4137 22276 4141 22332
rect 4077 22272 4141 22276
rect 4157 22332 4221 22336
rect 4157 22276 4161 22332
rect 4161 22276 4217 22332
rect 4217 22276 4221 22332
rect 4157 22272 4221 22276
rect 9848 22332 9912 22336
rect 9848 22276 9852 22332
rect 9852 22276 9908 22332
rect 9908 22276 9912 22332
rect 9848 22272 9912 22276
rect 9928 22332 9992 22336
rect 9928 22276 9932 22332
rect 9932 22276 9988 22332
rect 9988 22276 9992 22332
rect 9928 22272 9992 22276
rect 10008 22332 10072 22336
rect 10008 22276 10012 22332
rect 10012 22276 10068 22332
rect 10068 22276 10072 22332
rect 10008 22272 10072 22276
rect 10088 22332 10152 22336
rect 10088 22276 10092 22332
rect 10092 22276 10148 22332
rect 10148 22276 10152 22332
rect 10088 22272 10152 22276
rect 15778 22332 15842 22336
rect 15778 22276 15782 22332
rect 15782 22276 15838 22332
rect 15838 22276 15842 22332
rect 15778 22272 15842 22276
rect 15858 22332 15922 22336
rect 15858 22276 15862 22332
rect 15862 22276 15918 22332
rect 15918 22276 15922 22332
rect 15858 22272 15922 22276
rect 15938 22332 16002 22336
rect 15938 22276 15942 22332
rect 15942 22276 15998 22332
rect 15998 22276 16002 22332
rect 15938 22272 16002 22276
rect 16018 22332 16082 22336
rect 16018 22276 16022 22332
rect 16022 22276 16078 22332
rect 16078 22276 16082 22332
rect 16018 22272 16082 22276
rect 6882 21788 6946 21792
rect 6882 21732 6886 21788
rect 6886 21732 6942 21788
rect 6942 21732 6946 21788
rect 6882 21728 6946 21732
rect 6962 21788 7026 21792
rect 6962 21732 6966 21788
rect 6966 21732 7022 21788
rect 7022 21732 7026 21788
rect 6962 21728 7026 21732
rect 7042 21788 7106 21792
rect 7042 21732 7046 21788
rect 7046 21732 7102 21788
rect 7102 21732 7106 21788
rect 7042 21728 7106 21732
rect 7122 21788 7186 21792
rect 7122 21732 7126 21788
rect 7126 21732 7182 21788
rect 7182 21732 7186 21788
rect 7122 21728 7186 21732
rect 12813 21788 12877 21792
rect 12813 21732 12817 21788
rect 12817 21732 12873 21788
rect 12873 21732 12877 21788
rect 12813 21728 12877 21732
rect 12893 21788 12957 21792
rect 12893 21732 12897 21788
rect 12897 21732 12953 21788
rect 12953 21732 12957 21788
rect 12893 21728 12957 21732
rect 12973 21788 13037 21792
rect 12973 21732 12977 21788
rect 12977 21732 13033 21788
rect 13033 21732 13037 21788
rect 12973 21728 13037 21732
rect 13053 21788 13117 21792
rect 13053 21732 13057 21788
rect 13057 21732 13113 21788
rect 13113 21732 13117 21788
rect 13053 21728 13117 21732
rect 3917 21244 3981 21248
rect 3917 21188 3921 21244
rect 3921 21188 3977 21244
rect 3977 21188 3981 21244
rect 3917 21184 3981 21188
rect 3997 21244 4061 21248
rect 3997 21188 4001 21244
rect 4001 21188 4057 21244
rect 4057 21188 4061 21244
rect 3997 21184 4061 21188
rect 4077 21244 4141 21248
rect 4077 21188 4081 21244
rect 4081 21188 4137 21244
rect 4137 21188 4141 21244
rect 4077 21184 4141 21188
rect 4157 21244 4221 21248
rect 4157 21188 4161 21244
rect 4161 21188 4217 21244
rect 4217 21188 4221 21244
rect 4157 21184 4221 21188
rect 9848 21244 9912 21248
rect 9848 21188 9852 21244
rect 9852 21188 9908 21244
rect 9908 21188 9912 21244
rect 9848 21184 9912 21188
rect 9928 21244 9992 21248
rect 9928 21188 9932 21244
rect 9932 21188 9988 21244
rect 9988 21188 9992 21244
rect 9928 21184 9992 21188
rect 10008 21244 10072 21248
rect 10008 21188 10012 21244
rect 10012 21188 10068 21244
rect 10068 21188 10072 21244
rect 10008 21184 10072 21188
rect 10088 21244 10152 21248
rect 10088 21188 10092 21244
rect 10092 21188 10148 21244
rect 10148 21188 10152 21244
rect 10088 21184 10152 21188
rect 15778 21244 15842 21248
rect 15778 21188 15782 21244
rect 15782 21188 15838 21244
rect 15838 21188 15842 21244
rect 15778 21184 15842 21188
rect 15858 21244 15922 21248
rect 15858 21188 15862 21244
rect 15862 21188 15918 21244
rect 15918 21188 15922 21244
rect 15858 21184 15922 21188
rect 15938 21244 16002 21248
rect 15938 21188 15942 21244
rect 15942 21188 15998 21244
rect 15998 21188 16002 21244
rect 15938 21184 16002 21188
rect 16018 21244 16082 21248
rect 16018 21188 16022 21244
rect 16022 21188 16078 21244
rect 16078 21188 16082 21244
rect 16018 21184 16082 21188
rect 6882 20700 6946 20704
rect 6882 20644 6886 20700
rect 6886 20644 6942 20700
rect 6942 20644 6946 20700
rect 6882 20640 6946 20644
rect 6962 20700 7026 20704
rect 6962 20644 6966 20700
rect 6966 20644 7022 20700
rect 7022 20644 7026 20700
rect 6962 20640 7026 20644
rect 7042 20700 7106 20704
rect 7042 20644 7046 20700
rect 7046 20644 7102 20700
rect 7102 20644 7106 20700
rect 7042 20640 7106 20644
rect 7122 20700 7186 20704
rect 7122 20644 7126 20700
rect 7126 20644 7182 20700
rect 7182 20644 7186 20700
rect 7122 20640 7186 20644
rect 12813 20700 12877 20704
rect 12813 20644 12817 20700
rect 12817 20644 12873 20700
rect 12873 20644 12877 20700
rect 12813 20640 12877 20644
rect 12893 20700 12957 20704
rect 12893 20644 12897 20700
rect 12897 20644 12953 20700
rect 12953 20644 12957 20700
rect 12893 20640 12957 20644
rect 12973 20700 13037 20704
rect 12973 20644 12977 20700
rect 12977 20644 13033 20700
rect 13033 20644 13037 20700
rect 12973 20640 13037 20644
rect 13053 20700 13117 20704
rect 13053 20644 13057 20700
rect 13057 20644 13113 20700
rect 13113 20644 13117 20700
rect 13053 20640 13117 20644
rect 3917 20156 3981 20160
rect 3917 20100 3921 20156
rect 3921 20100 3977 20156
rect 3977 20100 3981 20156
rect 3917 20096 3981 20100
rect 3997 20156 4061 20160
rect 3997 20100 4001 20156
rect 4001 20100 4057 20156
rect 4057 20100 4061 20156
rect 3997 20096 4061 20100
rect 4077 20156 4141 20160
rect 4077 20100 4081 20156
rect 4081 20100 4137 20156
rect 4137 20100 4141 20156
rect 4077 20096 4141 20100
rect 4157 20156 4221 20160
rect 4157 20100 4161 20156
rect 4161 20100 4217 20156
rect 4217 20100 4221 20156
rect 4157 20096 4221 20100
rect 9848 20156 9912 20160
rect 9848 20100 9852 20156
rect 9852 20100 9908 20156
rect 9908 20100 9912 20156
rect 9848 20096 9912 20100
rect 9928 20156 9992 20160
rect 9928 20100 9932 20156
rect 9932 20100 9988 20156
rect 9988 20100 9992 20156
rect 9928 20096 9992 20100
rect 10008 20156 10072 20160
rect 10008 20100 10012 20156
rect 10012 20100 10068 20156
rect 10068 20100 10072 20156
rect 10008 20096 10072 20100
rect 10088 20156 10152 20160
rect 10088 20100 10092 20156
rect 10092 20100 10148 20156
rect 10148 20100 10152 20156
rect 10088 20096 10152 20100
rect 15778 20156 15842 20160
rect 15778 20100 15782 20156
rect 15782 20100 15838 20156
rect 15838 20100 15842 20156
rect 15778 20096 15842 20100
rect 15858 20156 15922 20160
rect 15858 20100 15862 20156
rect 15862 20100 15918 20156
rect 15918 20100 15922 20156
rect 15858 20096 15922 20100
rect 15938 20156 16002 20160
rect 15938 20100 15942 20156
rect 15942 20100 15998 20156
rect 15998 20100 16002 20156
rect 15938 20096 16002 20100
rect 16018 20156 16082 20160
rect 16018 20100 16022 20156
rect 16022 20100 16078 20156
rect 16078 20100 16082 20156
rect 16018 20096 16082 20100
rect 6882 19612 6946 19616
rect 6882 19556 6886 19612
rect 6886 19556 6942 19612
rect 6942 19556 6946 19612
rect 6882 19552 6946 19556
rect 6962 19612 7026 19616
rect 6962 19556 6966 19612
rect 6966 19556 7022 19612
rect 7022 19556 7026 19612
rect 6962 19552 7026 19556
rect 7042 19612 7106 19616
rect 7042 19556 7046 19612
rect 7046 19556 7102 19612
rect 7102 19556 7106 19612
rect 7042 19552 7106 19556
rect 7122 19612 7186 19616
rect 7122 19556 7126 19612
rect 7126 19556 7182 19612
rect 7182 19556 7186 19612
rect 7122 19552 7186 19556
rect 12813 19612 12877 19616
rect 12813 19556 12817 19612
rect 12817 19556 12873 19612
rect 12873 19556 12877 19612
rect 12813 19552 12877 19556
rect 12893 19612 12957 19616
rect 12893 19556 12897 19612
rect 12897 19556 12953 19612
rect 12953 19556 12957 19612
rect 12893 19552 12957 19556
rect 12973 19612 13037 19616
rect 12973 19556 12977 19612
rect 12977 19556 13033 19612
rect 13033 19556 13037 19612
rect 12973 19552 13037 19556
rect 13053 19612 13117 19616
rect 13053 19556 13057 19612
rect 13057 19556 13113 19612
rect 13113 19556 13117 19612
rect 13053 19552 13117 19556
rect 3917 19068 3981 19072
rect 3917 19012 3921 19068
rect 3921 19012 3977 19068
rect 3977 19012 3981 19068
rect 3917 19008 3981 19012
rect 3997 19068 4061 19072
rect 3997 19012 4001 19068
rect 4001 19012 4057 19068
rect 4057 19012 4061 19068
rect 3997 19008 4061 19012
rect 4077 19068 4141 19072
rect 4077 19012 4081 19068
rect 4081 19012 4137 19068
rect 4137 19012 4141 19068
rect 4077 19008 4141 19012
rect 4157 19068 4221 19072
rect 4157 19012 4161 19068
rect 4161 19012 4217 19068
rect 4217 19012 4221 19068
rect 4157 19008 4221 19012
rect 9848 19068 9912 19072
rect 9848 19012 9852 19068
rect 9852 19012 9908 19068
rect 9908 19012 9912 19068
rect 9848 19008 9912 19012
rect 9928 19068 9992 19072
rect 9928 19012 9932 19068
rect 9932 19012 9988 19068
rect 9988 19012 9992 19068
rect 9928 19008 9992 19012
rect 10008 19068 10072 19072
rect 10008 19012 10012 19068
rect 10012 19012 10068 19068
rect 10068 19012 10072 19068
rect 10008 19008 10072 19012
rect 10088 19068 10152 19072
rect 10088 19012 10092 19068
rect 10092 19012 10148 19068
rect 10148 19012 10152 19068
rect 10088 19008 10152 19012
rect 15778 19068 15842 19072
rect 15778 19012 15782 19068
rect 15782 19012 15838 19068
rect 15838 19012 15842 19068
rect 15778 19008 15842 19012
rect 15858 19068 15922 19072
rect 15858 19012 15862 19068
rect 15862 19012 15918 19068
rect 15918 19012 15922 19068
rect 15858 19008 15922 19012
rect 15938 19068 16002 19072
rect 15938 19012 15942 19068
rect 15942 19012 15998 19068
rect 15998 19012 16002 19068
rect 15938 19008 16002 19012
rect 16018 19068 16082 19072
rect 16018 19012 16022 19068
rect 16022 19012 16078 19068
rect 16078 19012 16082 19068
rect 16018 19008 16082 19012
rect 6882 18524 6946 18528
rect 6882 18468 6886 18524
rect 6886 18468 6942 18524
rect 6942 18468 6946 18524
rect 6882 18464 6946 18468
rect 6962 18524 7026 18528
rect 6962 18468 6966 18524
rect 6966 18468 7022 18524
rect 7022 18468 7026 18524
rect 6962 18464 7026 18468
rect 7042 18524 7106 18528
rect 7042 18468 7046 18524
rect 7046 18468 7102 18524
rect 7102 18468 7106 18524
rect 7042 18464 7106 18468
rect 7122 18524 7186 18528
rect 7122 18468 7126 18524
rect 7126 18468 7182 18524
rect 7182 18468 7186 18524
rect 7122 18464 7186 18468
rect 12813 18524 12877 18528
rect 12813 18468 12817 18524
rect 12817 18468 12873 18524
rect 12873 18468 12877 18524
rect 12813 18464 12877 18468
rect 12893 18524 12957 18528
rect 12893 18468 12897 18524
rect 12897 18468 12953 18524
rect 12953 18468 12957 18524
rect 12893 18464 12957 18468
rect 12973 18524 13037 18528
rect 12973 18468 12977 18524
rect 12977 18468 13033 18524
rect 13033 18468 13037 18524
rect 12973 18464 13037 18468
rect 13053 18524 13117 18528
rect 13053 18468 13057 18524
rect 13057 18468 13113 18524
rect 13113 18468 13117 18524
rect 13053 18464 13117 18468
rect 3917 17980 3981 17984
rect 3917 17924 3921 17980
rect 3921 17924 3977 17980
rect 3977 17924 3981 17980
rect 3917 17920 3981 17924
rect 3997 17980 4061 17984
rect 3997 17924 4001 17980
rect 4001 17924 4057 17980
rect 4057 17924 4061 17980
rect 3997 17920 4061 17924
rect 4077 17980 4141 17984
rect 4077 17924 4081 17980
rect 4081 17924 4137 17980
rect 4137 17924 4141 17980
rect 4077 17920 4141 17924
rect 4157 17980 4221 17984
rect 4157 17924 4161 17980
rect 4161 17924 4217 17980
rect 4217 17924 4221 17980
rect 4157 17920 4221 17924
rect 9848 17980 9912 17984
rect 9848 17924 9852 17980
rect 9852 17924 9908 17980
rect 9908 17924 9912 17980
rect 9848 17920 9912 17924
rect 9928 17980 9992 17984
rect 9928 17924 9932 17980
rect 9932 17924 9988 17980
rect 9988 17924 9992 17980
rect 9928 17920 9992 17924
rect 10008 17980 10072 17984
rect 10008 17924 10012 17980
rect 10012 17924 10068 17980
rect 10068 17924 10072 17980
rect 10008 17920 10072 17924
rect 10088 17980 10152 17984
rect 10088 17924 10092 17980
rect 10092 17924 10148 17980
rect 10148 17924 10152 17980
rect 10088 17920 10152 17924
rect 15778 17980 15842 17984
rect 15778 17924 15782 17980
rect 15782 17924 15838 17980
rect 15838 17924 15842 17980
rect 15778 17920 15842 17924
rect 15858 17980 15922 17984
rect 15858 17924 15862 17980
rect 15862 17924 15918 17980
rect 15918 17924 15922 17980
rect 15858 17920 15922 17924
rect 15938 17980 16002 17984
rect 15938 17924 15942 17980
rect 15942 17924 15998 17980
rect 15998 17924 16002 17980
rect 15938 17920 16002 17924
rect 16018 17980 16082 17984
rect 16018 17924 16022 17980
rect 16022 17924 16078 17980
rect 16078 17924 16082 17980
rect 16018 17920 16082 17924
rect 6882 17436 6946 17440
rect 6882 17380 6886 17436
rect 6886 17380 6942 17436
rect 6942 17380 6946 17436
rect 6882 17376 6946 17380
rect 6962 17436 7026 17440
rect 6962 17380 6966 17436
rect 6966 17380 7022 17436
rect 7022 17380 7026 17436
rect 6962 17376 7026 17380
rect 7042 17436 7106 17440
rect 7042 17380 7046 17436
rect 7046 17380 7102 17436
rect 7102 17380 7106 17436
rect 7042 17376 7106 17380
rect 7122 17436 7186 17440
rect 7122 17380 7126 17436
rect 7126 17380 7182 17436
rect 7182 17380 7186 17436
rect 7122 17376 7186 17380
rect 12813 17436 12877 17440
rect 12813 17380 12817 17436
rect 12817 17380 12873 17436
rect 12873 17380 12877 17436
rect 12813 17376 12877 17380
rect 12893 17436 12957 17440
rect 12893 17380 12897 17436
rect 12897 17380 12953 17436
rect 12953 17380 12957 17436
rect 12893 17376 12957 17380
rect 12973 17436 13037 17440
rect 12973 17380 12977 17436
rect 12977 17380 13033 17436
rect 13033 17380 13037 17436
rect 12973 17376 13037 17380
rect 13053 17436 13117 17440
rect 13053 17380 13057 17436
rect 13057 17380 13113 17436
rect 13113 17380 13117 17436
rect 13053 17376 13117 17380
rect 3917 16892 3981 16896
rect 3917 16836 3921 16892
rect 3921 16836 3977 16892
rect 3977 16836 3981 16892
rect 3917 16832 3981 16836
rect 3997 16892 4061 16896
rect 3997 16836 4001 16892
rect 4001 16836 4057 16892
rect 4057 16836 4061 16892
rect 3997 16832 4061 16836
rect 4077 16892 4141 16896
rect 4077 16836 4081 16892
rect 4081 16836 4137 16892
rect 4137 16836 4141 16892
rect 4077 16832 4141 16836
rect 4157 16892 4221 16896
rect 4157 16836 4161 16892
rect 4161 16836 4217 16892
rect 4217 16836 4221 16892
rect 4157 16832 4221 16836
rect 9848 16892 9912 16896
rect 9848 16836 9852 16892
rect 9852 16836 9908 16892
rect 9908 16836 9912 16892
rect 9848 16832 9912 16836
rect 9928 16892 9992 16896
rect 9928 16836 9932 16892
rect 9932 16836 9988 16892
rect 9988 16836 9992 16892
rect 9928 16832 9992 16836
rect 10008 16892 10072 16896
rect 10008 16836 10012 16892
rect 10012 16836 10068 16892
rect 10068 16836 10072 16892
rect 10008 16832 10072 16836
rect 10088 16892 10152 16896
rect 10088 16836 10092 16892
rect 10092 16836 10148 16892
rect 10148 16836 10152 16892
rect 10088 16832 10152 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 15938 16892 16002 16896
rect 15938 16836 15942 16892
rect 15942 16836 15998 16892
rect 15998 16836 16002 16892
rect 15938 16832 16002 16836
rect 16018 16892 16082 16896
rect 16018 16836 16022 16892
rect 16022 16836 16078 16892
rect 16078 16836 16082 16892
rect 16018 16832 16082 16836
rect 6882 16348 6946 16352
rect 6882 16292 6886 16348
rect 6886 16292 6942 16348
rect 6942 16292 6946 16348
rect 6882 16288 6946 16292
rect 6962 16348 7026 16352
rect 6962 16292 6966 16348
rect 6966 16292 7022 16348
rect 7022 16292 7026 16348
rect 6962 16288 7026 16292
rect 7042 16348 7106 16352
rect 7042 16292 7046 16348
rect 7046 16292 7102 16348
rect 7102 16292 7106 16348
rect 7042 16288 7106 16292
rect 7122 16348 7186 16352
rect 7122 16292 7126 16348
rect 7126 16292 7182 16348
rect 7182 16292 7186 16348
rect 7122 16288 7186 16292
rect 12813 16348 12877 16352
rect 12813 16292 12817 16348
rect 12817 16292 12873 16348
rect 12873 16292 12877 16348
rect 12813 16288 12877 16292
rect 12893 16348 12957 16352
rect 12893 16292 12897 16348
rect 12897 16292 12953 16348
rect 12953 16292 12957 16348
rect 12893 16288 12957 16292
rect 12973 16348 13037 16352
rect 12973 16292 12977 16348
rect 12977 16292 13033 16348
rect 13033 16292 13037 16348
rect 12973 16288 13037 16292
rect 13053 16348 13117 16352
rect 13053 16292 13057 16348
rect 13057 16292 13113 16348
rect 13113 16292 13117 16348
rect 13053 16288 13117 16292
rect 3917 15804 3981 15808
rect 3917 15748 3921 15804
rect 3921 15748 3977 15804
rect 3977 15748 3981 15804
rect 3917 15744 3981 15748
rect 3997 15804 4061 15808
rect 3997 15748 4001 15804
rect 4001 15748 4057 15804
rect 4057 15748 4061 15804
rect 3997 15744 4061 15748
rect 4077 15804 4141 15808
rect 4077 15748 4081 15804
rect 4081 15748 4137 15804
rect 4137 15748 4141 15804
rect 4077 15744 4141 15748
rect 4157 15804 4221 15808
rect 4157 15748 4161 15804
rect 4161 15748 4217 15804
rect 4217 15748 4221 15804
rect 4157 15744 4221 15748
rect 9848 15804 9912 15808
rect 9848 15748 9852 15804
rect 9852 15748 9908 15804
rect 9908 15748 9912 15804
rect 9848 15744 9912 15748
rect 9928 15804 9992 15808
rect 9928 15748 9932 15804
rect 9932 15748 9988 15804
rect 9988 15748 9992 15804
rect 9928 15744 9992 15748
rect 10008 15804 10072 15808
rect 10008 15748 10012 15804
rect 10012 15748 10068 15804
rect 10068 15748 10072 15804
rect 10008 15744 10072 15748
rect 10088 15804 10152 15808
rect 10088 15748 10092 15804
rect 10092 15748 10148 15804
rect 10148 15748 10152 15804
rect 10088 15744 10152 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 15938 15804 16002 15808
rect 15938 15748 15942 15804
rect 15942 15748 15998 15804
rect 15998 15748 16002 15804
rect 15938 15744 16002 15748
rect 16018 15804 16082 15808
rect 16018 15748 16022 15804
rect 16022 15748 16078 15804
rect 16078 15748 16082 15804
rect 16018 15744 16082 15748
rect 6882 15260 6946 15264
rect 6882 15204 6886 15260
rect 6886 15204 6942 15260
rect 6942 15204 6946 15260
rect 6882 15200 6946 15204
rect 6962 15260 7026 15264
rect 6962 15204 6966 15260
rect 6966 15204 7022 15260
rect 7022 15204 7026 15260
rect 6962 15200 7026 15204
rect 7042 15260 7106 15264
rect 7042 15204 7046 15260
rect 7046 15204 7102 15260
rect 7102 15204 7106 15260
rect 7042 15200 7106 15204
rect 7122 15260 7186 15264
rect 7122 15204 7126 15260
rect 7126 15204 7182 15260
rect 7182 15204 7186 15260
rect 7122 15200 7186 15204
rect 12813 15260 12877 15264
rect 12813 15204 12817 15260
rect 12817 15204 12873 15260
rect 12873 15204 12877 15260
rect 12813 15200 12877 15204
rect 12893 15260 12957 15264
rect 12893 15204 12897 15260
rect 12897 15204 12953 15260
rect 12953 15204 12957 15260
rect 12893 15200 12957 15204
rect 12973 15260 13037 15264
rect 12973 15204 12977 15260
rect 12977 15204 13033 15260
rect 13033 15204 13037 15260
rect 12973 15200 13037 15204
rect 13053 15260 13117 15264
rect 13053 15204 13057 15260
rect 13057 15204 13113 15260
rect 13113 15204 13117 15260
rect 13053 15200 13117 15204
rect 3917 14716 3981 14720
rect 3917 14660 3921 14716
rect 3921 14660 3977 14716
rect 3977 14660 3981 14716
rect 3917 14656 3981 14660
rect 3997 14716 4061 14720
rect 3997 14660 4001 14716
rect 4001 14660 4057 14716
rect 4057 14660 4061 14716
rect 3997 14656 4061 14660
rect 4077 14716 4141 14720
rect 4077 14660 4081 14716
rect 4081 14660 4137 14716
rect 4137 14660 4141 14716
rect 4077 14656 4141 14660
rect 4157 14716 4221 14720
rect 4157 14660 4161 14716
rect 4161 14660 4217 14716
rect 4217 14660 4221 14716
rect 4157 14656 4221 14660
rect 9848 14716 9912 14720
rect 9848 14660 9852 14716
rect 9852 14660 9908 14716
rect 9908 14660 9912 14716
rect 9848 14656 9912 14660
rect 9928 14716 9992 14720
rect 9928 14660 9932 14716
rect 9932 14660 9988 14716
rect 9988 14660 9992 14716
rect 9928 14656 9992 14660
rect 10008 14716 10072 14720
rect 10008 14660 10012 14716
rect 10012 14660 10068 14716
rect 10068 14660 10072 14716
rect 10008 14656 10072 14660
rect 10088 14716 10152 14720
rect 10088 14660 10092 14716
rect 10092 14660 10148 14716
rect 10148 14660 10152 14716
rect 10088 14656 10152 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 15938 14716 16002 14720
rect 15938 14660 15942 14716
rect 15942 14660 15998 14716
rect 15998 14660 16002 14716
rect 15938 14656 16002 14660
rect 16018 14716 16082 14720
rect 16018 14660 16022 14716
rect 16022 14660 16078 14716
rect 16078 14660 16082 14716
rect 16018 14656 16082 14660
rect 6882 14172 6946 14176
rect 6882 14116 6886 14172
rect 6886 14116 6942 14172
rect 6942 14116 6946 14172
rect 6882 14112 6946 14116
rect 6962 14172 7026 14176
rect 6962 14116 6966 14172
rect 6966 14116 7022 14172
rect 7022 14116 7026 14172
rect 6962 14112 7026 14116
rect 7042 14172 7106 14176
rect 7042 14116 7046 14172
rect 7046 14116 7102 14172
rect 7102 14116 7106 14172
rect 7042 14112 7106 14116
rect 7122 14172 7186 14176
rect 7122 14116 7126 14172
rect 7126 14116 7182 14172
rect 7182 14116 7186 14172
rect 7122 14112 7186 14116
rect 12813 14172 12877 14176
rect 12813 14116 12817 14172
rect 12817 14116 12873 14172
rect 12873 14116 12877 14172
rect 12813 14112 12877 14116
rect 12893 14172 12957 14176
rect 12893 14116 12897 14172
rect 12897 14116 12953 14172
rect 12953 14116 12957 14172
rect 12893 14112 12957 14116
rect 12973 14172 13037 14176
rect 12973 14116 12977 14172
rect 12977 14116 13033 14172
rect 13033 14116 13037 14172
rect 12973 14112 13037 14116
rect 13053 14172 13117 14176
rect 13053 14116 13057 14172
rect 13057 14116 13113 14172
rect 13113 14116 13117 14172
rect 13053 14112 13117 14116
rect 3917 13628 3981 13632
rect 3917 13572 3921 13628
rect 3921 13572 3977 13628
rect 3977 13572 3981 13628
rect 3917 13568 3981 13572
rect 3997 13628 4061 13632
rect 3997 13572 4001 13628
rect 4001 13572 4057 13628
rect 4057 13572 4061 13628
rect 3997 13568 4061 13572
rect 4077 13628 4141 13632
rect 4077 13572 4081 13628
rect 4081 13572 4137 13628
rect 4137 13572 4141 13628
rect 4077 13568 4141 13572
rect 4157 13628 4221 13632
rect 4157 13572 4161 13628
rect 4161 13572 4217 13628
rect 4217 13572 4221 13628
rect 4157 13568 4221 13572
rect 9848 13628 9912 13632
rect 9848 13572 9852 13628
rect 9852 13572 9908 13628
rect 9908 13572 9912 13628
rect 9848 13568 9912 13572
rect 9928 13628 9992 13632
rect 9928 13572 9932 13628
rect 9932 13572 9988 13628
rect 9988 13572 9992 13628
rect 9928 13568 9992 13572
rect 10008 13628 10072 13632
rect 10008 13572 10012 13628
rect 10012 13572 10068 13628
rect 10068 13572 10072 13628
rect 10008 13568 10072 13572
rect 10088 13628 10152 13632
rect 10088 13572 10092 13628
rect 10092 13572 10148 13628
rect 10148 13572 10152 13628
rect 10088 13568 10152 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 15938 13628 16002 13632
rect 15938 13572 15942 13628
rect 15942 13572 15998 13628
rect 15998 13572 16002 13628
rect 15938 13568 16002 13572
rect 16018 13628 16082 13632
rect 16018 13572 16022 13628
rect 16022 13572 16078 13628
rect 16078 13572 16082 13628
rect 16018 13568 16082 13572
rect 6882 13084 6946 13088
rect 6882 13028 6886 13084
rect 6886 13028 6942 13084
rect 6942 13028 6946 13084
rect 6882 13024 6946 13028
rect 6962 13084 7026 13088
rect 6962 13028 6966 13084
rect 6966 13028 7022 13084
rect 7022 13028 7026 13084
rect 6962 13024 7026 13028
rect 7042 13084 7106 13088
rect 7042 13028 7046 13084
rect 7046 13028 7102 13084
rect 7102 13028 7106 13084
rect 7042 13024 7106 13028
rect 7122 13084 7186 13088
rect 7122 13028 7126 13084
rect 7126 13028 7182 13084
rect 7182 13028 7186 13084
rect 7122 13024 7186 13028
rect 12813 13084 12877 13088
rect 12813 13028 12817 13084
rect 12817 13028 12873 13084
rect 12873 13028 12877 13084
rect 12813 13024 12877 13028
rect 12893 13084 12957 13088
rect 12893 13028 12897 13084
rect 12897 13028 12953 13084
rect 12953 13028 12957 13084
rect 12893 13024 12957 13028
rect 12973 13084 13037 13088
rect 12973 13028 12977 13084
rect 12977 13028 13033 13084
rect 13033 13028 13037 13084
rect 12973 13024 13037 13028
rect 13053 13084 13117 13088
rect 13053 13028 13057 13084
rect 13057 13028 13113 13084
rect 13113 13028 13117 13084
rect 13053 13024 13117 13028
rect 3917 12540 3981 12544
rect 3917 12484 3921 12540
rect 3921 12484 3977 12540
rect 3977 12484 3981 12540
rect 3917 12480 3981 12484
rect 3997 12540 4061 12544
rect 3997 12484 4001 12540
rect 4001 12484 4057 12540
rect 4057 12484 4061 12540
rect 3997 12480 4061 12484
rect 4077 12540 4141 12544
rect 4077 12484 4081 12540
rect 4081 12484 4137 12540
rect 4137 12484 4141 12540
rect 4077 12480 4141 12484
rect 4157 12540 4221 12544
rect 4157 12484 4161 12540
rect 4161 12484 4217 12540
rect 4217 12484 4221 12540
rect 4157 12480 4221 12484
rect 9848 12540 9912 12544
rect 9848 12484 9852 12540
rect 9852 12484 9908 12540
rect 9908 12484 9912 12540
rect 9848 12480 9912 12484
rect 9928 12540 9992 12544
rect 9928 12484 9932 12540
rect 9932 12484 9988 12540
rect 9988 12484 9992 12540
rect 9928 12480 9992 12484
rect 10008 12540 10072 12544
rect 10008 12484 10012 12540
rect 10012 12484 10068 12540
rect 10068 12484 10072 12540
rect 10008 12480 10072 12484
rect 10088 12540 10152 12544
rect 10088 12484 10092 12540
rect 10092 12484 10148 12540
rect 10148 12484 10152 12540
rect 10088 12480 10152 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 15938 12540 16002 12544
rect 15938 12484 15942 12540
rect 15942 12484 15998 12540
rect 15998 12484 16002 12540
rect 15938 12480 16002 12484
rect 16018 12540 16082 12544
rect 16018 12484 16022 12540
rect 16022 12484 16078 12540
rect 16078 12484 16082 12540
rect 16018 12480 16082 12484
rect 6882 11996 6946 12000
rect 6882 11940 6886 11996
rect 6886 11940 6942 11996
rect 6942 11940 6946 11996
rect 6882 11936 6946 11940
rect 6962 11996 7026 12000
rect 6962 11940 6966 11996
rect 6966 11940 7022 11996
rect 7022 11940 7026 11996
rect 6962 11936 7026 11940
rect 7042 11996 7106 12000
rect 7042 11940 7046 11996
rect 7046 11940 7102 11996
rect 7102 11940 7106 11996
rect 7042 11936 7106 11940
rect 7122 11996 7186 12000
rect 7122 11940 7126 11996
rect 7126 11940 7182 11996
rect 7182 11940 7186 11996
rect 7122 11936 7186 11940
rect 12813 11996 12877 12000
rect 12813 11940 12817 11996
rect 12817 11940 12873 11996
rect 12873 11940 12877 11996
rect 12813 11936 12877 11940
rect 12893 11996 12957 12000
rect 12893 11940 12897 11996
rect 12897 11940 12953 11996
rect 12953 11940 12957 11996
rect 12893 11936 12957 11940
rect 12973 11996 13037 12000
rect 12973 11940 12977 11996
rect 12977 11940 13033 11996
rect 13033 11940 13037 11996
rect 12973 11936 13037 11940
rect 13053 11996 13117 12000
rect 13053 11940 13057 11996
rect 13057 11940 13113 11996
rect 13113 11940 13117 11996
rect 13053 11936 13117 11940
rect 3917 11452 3981 11456
rect 3917 11396 3921 11452
rect 3921 11396 3977 11452
rect 3977 11396 3981 11452
rect 3917 11392 3981 11396
rect 3997 11452 4061 11456
rect 3997 11396 4001 11452
rect 4001 11396 4057 11452
rect 4057 11396 4061 11452
rect 3997 11392 4061 11396
rect 4077 11452 4141 11456
rect 4077 11396 4081 11452
rect 4081 11396 4137 11452
rect 4137 11396 4141 11452
rect 4077 11392 4141 11396
rect 4157 11452 4221 11456
rect 4157 11396 4161 11452
rect 4161 11396 4217 11452
rect 4217 11396 4221 11452
rect 4157 11392 4221 11396
rect 9848 11452 9912 11456
rect 9848 11396 9852 11452
rect 9852 11396 9908 11452
rect 9908 11396 9912 11452
rect 9848 11392 9912 11396
rect 9928 11452 9992 11456
rect 9928 11396 9932 11452
rect 9932 11396 9988 11452
rect 9988 11396 9992 11452
rect 9928 11392 9992 11396
rect 10008 11452 10072 11456
rect 10008 11396 10012 11452
rect 10012 11396 10068 11452
rect 10068 11396 10072 11452
rect 10008 11392 10072 11396
rect 10088 11452 10152 11456
rect 10088 11396 10092 11452
rect 10092 11396 10148 11452
rect 10148 11396 10152 11452
rect 10088 11392 10152 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 15938 11452 16002 11456
rect 15938 11396 15942 11452
rect 15942 11396 15998 11452
rect 15998 11396 16002 11452
rect 15938 11392 16002 11396
rect 16018 11452 16082 11456
rect 16018 11396 16022 11452
rect 16022 11396 16078 11452
rect 16078 11396 16082 11452
rect 16018 11392 16082 11396
rect 6882 10908 6946 10912
rect 6882 10852 6886 10908
rect 6886 10852 6942 10908
rect 6942 10852 6946 10908
rect 6882 10848 6946 10852
rect 6962 10908 7026 10912
rect 6962 10852 6966 10908
rect 6966 10852 7022 10908
rect 7022 10852 7026 10908
rect 6962 10848 7026 10852
rect 7042 10908 7106 10912
rect 7042 10852 7046 10908
rect 7046 10852 7102 10908
rect 7102 10852 7106 10908
rect 7042 10848 7106 10852
rect 7122 10908 7186 10912
rect 7122 10852 7126 10908
rect 7126 10852 7182 10908
rect 7182 10852 7186 10908
rect 7122 10848 7186 10852
rect 12813 10908 12877 10912
rect 12813 10852 12817 10908
rect 12817 10852 12873 10908
rect 12873 10852 12877 10908
rect 12813 10848 12877 10852
rect 12893 10908 12957 10912
rect 12893 10852 12897 10908
rect 12897 10852 12953 10908
rect 12953 10852 12957 10908
rect 12893 10848 12957 10852
rect 12973 10908 13037 10912
rect 12973 10852 12977 10908
rect 12977 10852 13033 10908
rect 13033 10852 13037 10908
rect 12973 10848 13037 10852
rect 13053 10908 13117 10912
rect 13053 10852 13057 10908
rect 13057 10852 13113 10908
rect 13113 10852 13117 10908
rect 13053 10848 13117 10852
rect 3917 10364 3981 10368
rect 3917 10308 3921 10364
rect 3921 10308 3977 10364
rect 3977 10308 3981 10364
rect 3917 10304 3981 10308
rect 3997 10364 4061 10368
rect 3997 10308 4001 10364
rect 4001 10308 4057 10364
rect 4057 10308 4061 10364
rect 3997 10304 4061 10308
rect 4077 10364 4141 10368
rect 4077 10308 4081 10364
rect 4081 10308 4137 10364
rect 4137 10308 4141 10364
rect 4077 10304 4141 10308
rect 4157 10364 4221 10368
rect 4157 10308 4161 10364
rect 4161 10308 4217 10364
rect 4217 10308 4221 10364
rect 4157 10304 4221 10308
rect 9848 10364 9912 10368
rect 9848 10308 9852 10364
rect 9852 10308 9908 10364
rect 9908 10308 9912 10364
rect 9848 10304 9912 10308
rect 9928 10364 9992 10368
rect 9928 10308 9932 10364
rect 9932 10308 9988 10364
rect 9988 10308 9992 10364
rect 9928 10304 9992 10308
rect 10008 10364 10072 10368
rect 10008 10308 10012 10364
rect 10012 10308 10068 10364
rect 10068 10308 10072 10364
rect 10008 10304 10072 10308
rect 10088 10364 10152 10368
rect 10088 10308 10092 10364
rect 10092 10308 10148 10364
rect 10148 10308 10152 10364
rect 10088 10304 10152 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 15938 10364 16002 10368
rect 15938 10308 15942 10364
rect 15942 10308 15998 10364
rect 15998 10308 16002 10364
rect 15938 10304 16002 10308
rect 16018 10364 16082 10368
rect 16018 10308 16022 10364
rect 16022 10308 16078 10364
rect 16078 10308 16082 10364
rect 16018 10304 16082 10308
rect 6882 9820 6946 9824
rect 6882 9764 6886 9820
rect 6886 9764 6942 9820
rect 6942 9764 6946 9820
rect 6882 9760 6946 9764
rect 6962 9820 7026 9824
rect 6962 9764 6966 9820
rect 6966 9764 7022 9820
rect 7022 9764 7026 9820
rect 6962 9760 7026 9764
rect 7042 9820 7106 9824
rect 7042 9764 7046 9820
rect 7046 9764 7102 9820
rect 7102 9764 7106 9820
rect 7042 9760 7106 9764
rect 7122 9820 7186 9824
rect 7122 9764 7126 9820
rect 7126 9764 7182 9820
rect 7182 9764 7186 9820
rect 7122 9760 7186 9764
rect 12813 9820 12877 9824
rect 12813 9764 12817 9820
rect 12817 9764 12873 9820
rect 12873 9764 12877 9820
rect 12813 9760 12877 9764
rect 12893 9820 12957 9824
rect 12893 9764 12897 9820
rect 12897 9764 12953 9820
rect 12953 9764 12957 9820
rect 12893 9760 12957 9764
rect 12973 9820 13037 9824
rect 12973 9764 12977 9820
rect 12977 9764 13033 9820
rect 13033 9764 13037 9820
rect 12973 9760 13037 9764
rect 13053 9820 13117 9824
rect 13053 9764 13057 9820
rect 13057 9764 13113 9820
rect 13113 9764 13117 9820
rect 13053 9760 13117 9764
rect 3917 9276 3981 9280
rect 3917 9220 3921 9276
rect 3921 9220 3977 9276
rect 3977 9220 3981 9276
rect 3917 9216 3981 9220
rect 3997 9276 4061 9280
rect 3997 9220 4001 9276
rect 4001 9220 4057 9276
rect 4057 9220 4061 9276
rect 3997 9216 4061 9220
rect 4077 9276 4141 9280
rect 4077 9220 4081 9276
rect 4081 9220 4137 9276
rect 4137 9220 4141 9276
rect 4077 9216 4141 9220
rect 4157 9276 4221 9280
rect 4157 9220 4161 9276
rect 4161 9220 4217 9276
rect 4217 9220 4221 9276
rect 4157 9216 4221 9220
rect 9848 9276 9912 9280
rect 9848 9220 9852 9276
rect 9852 9220 9908 9276
rect 9908 9220 9912 9276
rect 9848 9216 9912 9220
rect 9928 9276 9992 9280
rect 9928 9220 9932 9276
rect 9932 9220 9988 9276
rect 9988 9220 9992 9276
rect 9928 9216 9992 9220
rect 10008 9276 10072 9280
rect 10008 9220 10012 9276
rect 10012 9220 10068 9276
rect 10068 9220 10072 9276
rect 10008 9216 10072 9220
rect 10088 9276 10152 9280
rect 10088 9220 10092 9276
rect 10092 9220 10148 9276
rect 10148 9220 10152 9276
rect 10088 9216 10152 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 15938 9276 16002 9280
rect 15938 9220 15942 9276
rect 15942 9220 15998 9276
rect 15998 9220 16002 9276
rect 15938 9216 16002 9220
rect 16018 9276 16082 9280
rect 16018 9220 16022 9276
rect 16022 9220 16078 9276
rect 16078 9220 16082 9276
rect 16018 9216 16082 9220
rect 6882 8732 6946 8736
rect 6882 8676 6886 8732
rect 6886 8676 6942 8732
rect 6942 8676 6946 8732
rect 6882 8672 6946 8676
rect 6962 8732 7026 8736
rect 6962 8676 6966 8732
rect 6966 8676 7022 8732
rect 7022 8676 7026 8732
rect 6962 8672 7026 8676
rect 7042 8732 7106 8736
rect 7042 8676 7046 8732
rect 7046 8676 7102 8732
rect 7102 8676 7106 8732
rect 7042 8672 7106 8676
rect 7122 8732 7186 8736
rect 7122 8676 7126 8732
rect 7126 8676 7182 8732
rect 7182 8676 7186 8732
rect 7122 8672 7186 8676
rect 12813 8732 12877 8736
rect 12813 8676 12817 8732
rect 12817 8676 12873 8732
rect 12873 8676 12877 8732
rect 12813 8672 12877 8676
rect 12893 8732 12957 8736
rect 12893 8676 12897 8732
rect 12897 8676 12953 8732
rect 12953 8676 12957 8732
rect 12893 8672 12957 8676
rect 12973 8732 13037 8736
rect 12973 8676 12977 8732
rect 12977 8676 13033 8732
rect 13033 8676 13037 8732
rect 12973 8672 13037 8676
rect 13053 8732 13117 8736
rect 13053 8676 13057 8732
rect 13057 8676 13113 8732
rect 13113 8676 13117 8732
rect 13053 8672 13117 8676
rect 3917 8188 3981 8192
rect 3917 8132 3921 8188
rect 3921 8132 3977 8188
rect 3977 8132 3981 8188
rect 3917 8128 3981 8132
rect 3997 8188 4061 8192
rect 3997 8132 4001 8188
rect 4001 8132 4057 8188
rect 4057 8132 4061 8188
rect 3997 8128 4061 8132
rect 4077 8188 4141 8192
rect 4077 8132 4081 8188
rect 4081 8132 4137 8188
rect 4137 8132 4141 8188
rect 4077 8128 4141 8132
rect 4157 8188 4221 8192
rect 4157 8132 4161 8188
rect 4161 8132 4217 8188
rect 4217 8132 4221 8188
rect 4157 8128 4221 8132
rect 9848 8188 9912 8192
rect 9848 8132 9852 8188
rect 9852 8132 9908 8188
rect 9908 8132 9912 8188
rect 9848 8128 9912 8132
rect 9928 8188 9992 8192
rect 9928 8132 9932 8188
rect 9932 8132 9988 8188
rect 9988 8132 9992 8188
rect 9928 8128 9992 8132
rect 10008 8188 10072 8192
rect 10008 8132 10012 8188
rect 10012 8132 10068 8188
rect 10068 8132 10072 8188
rect 10008 8128 10072 8132
rect 10088 8188 10152 8192
rect 10088 8132 10092 8188
rect 10092 8132 10148 8188
rect 10148 8132 10152 8188
rect 10088 8128 10152 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 15938 8188 16002 8192
rect 15938 8132 15942 8188
rect 15942 8132 15998 8188
rect 15998 8132 16002 8188
rect 15938 8128 16002 8132
rect 16018 8188 16082 8192
rect 16018 8132 16022 8188
rect 16022 8132 16078 8188
rect 16078 8132 16082 8188
rect 16018 8128 16082 8132
rect 6882 7644 6946 7648
rect 6882 7588 6886 7644
rect 6886 7588 6942 7644
rect 6942 7588 6946 7644
rect 6882 7584 6946 7588
rect 6962 7644 7026 7648
rect 6962 7588 6966 7644
rect 6966 7588 7022 7644
rect 7022 7588 7026 7644
rect 6962 7584 7026 7588
rect 7042 7644 7106 7648
rect 7042 7588 7046 7644
rect 7046 7588 7102 7644
rect 7102 7588 7106 7644
rect 7042 7584 7106 7588
rect 7122 7644 7186 7648
rect 7122 7588 7126 7644
rect 7126 7588 7182 7644
rect 7182 7588 7186 7644
rect 7122 7584 7186 7588
rect 12813 7644 12877 7648
rect 12813 7588 12817 7644
rect 12817 7588 12873 7644
rect 12873 7588 12877 7644
rect 12813 7584 12877 7588
rect 12893 7644 12957 7648
rect 12893 7588 12897 7644
rect 12897 7588 12953 7644
rect 12953 7588 12957 7644
rect 12893 7584 12957 7588
rect 12973 7644 13037 7648
rect 12973 7588 12977 7644
rect 12977 7588 13033 7644
rect 13033 7588 13037 7644
rect 12973 7584 13037 7588
rect 13053 7644 13117 7648
rect 13053 7588 13057 7644
rect 13057 7588 13113 7644
rect 13113 7588 13117 7644
rect 13053 7584 13117 7588
rect 3917 7100 3981 7104
rect 3917 7044 3921 7100
rect 3921 7044 3977 7100
rect 3977 7044 3981 7100
rect 3917 7040 3981 7044
rect 3997 7100 4061 7104
rect 3997 7044 4001 7100
rect 4001 7044 4057 7100
rect 4057 7044 4061 7100
rect 3997 7040 4061 7044
rect 4077 7100 4141 7104
rect 4077 7044 4081 7100
rect 4081 7044 4137 7100
rect 4137 7044 4141 7100
rect 4077 7040 4141 7044
rect 4157 7100 4221 7104
rect 4157 7044 4161 7100
rect 4161 7044 4217 7100
rect 4217 7044 4221 7100
rect 4157 7040 4221 7044
rect 9848 7100 9912 7104
rect 9848 7044 9852 7100
rect 9852 7044 9908 7100
rect 9908 7044 9912 7100
rect 9848 7040 9912 7044
rect 9928 7100 9992 7104
rect 9928 7044 9932 7100
rect 9932 7044 9988 7100
rect 9988 7044 9992 7100
rect 9928 7040 9992 7044
rect 10008 7100 10072 7104
rect 10008 7044 10012 7100
rect 10012 7044 10068 7100
rect 10068 7044 10072 7100
rect 10008 7040 10072 7044
rect 10088 7100 10152 7104
rect 10088 7044 10092 7100
rect 10092 7044 10148 7100
rect 10148 7044 10152 7100
rect 10088 7040 10152 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 15938 7100 16002 7104
rect 15938 7044 15942 7100
rect 15942 7044 15998 7100
rect 15998 7044 16002 7100
rect 15938 7040 16002 7044
rect 16018 7100 16082 7104
rect 16018 7044 16022 7100
rect 16022 7044 16078 7100
rect 16078 7044 16082 7100
rect 16018 7040 16082 7044
rect 6882 6556 6946 6560
rect 6882 6500 6886 6556
rect 6886 6500 6942 6556
rect 6942 6500 6946 6556
rect 6882 6496 6946 6500
rect 6962 6556 7026 6560
rect 6962 6500 6966 6556
rect 6966 6500 7022 6556
rect 7022 6500 7026 6556
rect 6962 6496 7026 6500
rect 7042 6556 7106 6560
rect 7042 6500 7046 6556
rect 7046 6500 7102 6556
rect 7102 6500 7106 6556
rect 7042 6496 7106 6500
rect 7122 6556 7186 6560
rect 7122 6500 7126 6556
rect 7126 6500 7182 6556
rect 7182 6500 7186 6556
rect 7122 6496 7186 6500
rect 12813 6556 12877 6560
rect 12813 6500 12817 6556
rect 12817 6500 12873 6556
rect 12873 6500 12877 6556
rect 12813 6496 12877 6500
rect 12893 6556 12957 6560
rect 12893 6500 12897 6556
rect 12897 6500 12953 6556
rect 12953 6500 12957 6556
rect 12893 6496 12957 6500
rect 12973 6556 13037 6560
rect 12973 6500 12977 6556
rect 12977 6500 13033 6556
rect 13033 6500 13037 6556
rect 12973 6496 13037 6500
rect 13053 6556 13117 6560
rect 13053 6500 13057 6556
rect 13057 6500 13113 6556
rect 13113 6500 13117 6556
rect 13053 6496 13117 6500
rect 3917 6012 3981 6016
rect 3917 5956 3921 6012
rect 3921 5956 3977 6012
rect 3977 5956 3981 6012
rect 3917 5952 3981 5956
rect 3997 6012 4061 6016
rect 3997 5956 4001 6012
rect 4001 5956 4057 6012
rect 4057 5956 4061 6012
rect 3997 5952 4061 5956
rect 4077 6012 4141 6016
rect 4077 5956 4081 6012
rect 4081 5956 4137 6012
rect 4137 5956 4141 6012
rect 4077 5952 4141 5956
rect 4157 6012 4221 6016
rect 4157 5956 4161 6012
rect 4161 5956 4217 6012
rect 4217 5956 4221 6012
rect 4157 5952 4221 5956
rect 9848 6012 9912 6016
rect 9848 5956 9852 6012
rect 9852 5956 9908 6012
rect 9908 5956 9912 6012
rect 9848 5952 9912 5956
rect 9928 6012 9992 6016
rect 9928 5956 9932 6012
rect 9932 5956 9988 6012
rect 9988 5956 9992 6012
rect 9928 5952 9992 5956
rect 10008 6012 10072 6016
rect 10008 5956 10012 6012
rect 10012 5956 10068 6012
rect 10068 5956 10072 6012
rect 10008 5952 10072 5956
rect 10088 6012 10152 6016
rect 10088 5956 10092 6012
rect 10092 5956 10148 6012
rect 10148 5956 10152 6012
rect 10088 5952 10152 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 15938 6012 16002 6016
rect 15938 5956 15942 6012
rect 15942 5956 15998 6012
rect 15998 5956 16002 6012
rect 15938 5952 16002 5956
rect 16018 6012 16082 6016
rect 16018 5956 16022 6012
rect 16022 5956 16078 6012
rect 16078 5956 16082 6012
rect 16018 5952 16082 5956
rect 6882 5468 6946 5472
rect 6882 5412 6886 5468
rect 6886 5412 6942 5468
rect 6942 5412 6946 5468
rect 6882 5408 6946 5412
rect 6962 5468 7026 5472
rect 6962 5412 6966 5468
rect 6966 5412 7022 5468
rect 7022 5412 7026 5468
rect 6962 5408 7026 5412
rect 7042 5468 7106 5472
rect 7042 5412 7046 5468
rect 7046 5412 7102 5468
rect 7102 5412 7106 5468
rect 7042 5408 7106 5412
rect 7122 5468 7186 5472
rect 7122 5412 7126 5468
rect 7126 5412 7182 5468
rect 7182 5412 7186 5468
rect 7122 5408 7186 5412
rect 12813 5468 12877 5472
rect 12813 5412 12817 5468
rect 12817 5412 12873 5468
rect 12873 5412 12877 5468
rect 12813 5408 12877 5412
rect 12893 5468 12957 5472
rect 12893 5412 12897 5468
rect 12897 5412 12953 5468
rect 12953 5412 12957 5468
rect 12893 5408 12957 5412
rect 12973 5468 13037 5472
rect 12973 5412 12977 5468
rect 12977 5412 13033 5468
rect 13033 5412 13037 5468
rect 12973 5408 13037 5412
rect 13053 5468 13117 5472
rect 13053 5412 13057 5468
rect 13057 5412 13113 5468
rect 13113 5412 13117 5468
rect 13053 5408 13117 5412
rect 3917 4924 3981 4928
rect 3917 4868 3921 4924
rect 3921 4868 3977 4924
rect 3977 4868 3981 4924
rect 3917 4864 3981 4868
rect 3997 4924 4061 4928
rect 3997 4868 4001 4924
rect 4001 4868 4057 4924
rect 4057 4868 4061 4924
rect 3997 4864 4061 4868
rect 4077 4924 4141 4928
rect 4077 4868 4081 4924
rect 4081 4868 4137 4924
rect 4137 4868 4141 4924
rect 4077 4864 4141 4868
rect 4157 4924 4221 4928
rect 4157 4868 4161 4924
rect 4161 4868 4217 4924
rect 4217 4868 4221 4924
rect 4157 4864 4221 4868
rect 9848 4924 9912 4928
rect 9848 4868 9852 4924
rect 9852 4868 9908 4924
rect 9908 4868 9912 4924
rect 9848 4864 9912 4868
rect 9928 4924 9992 4928
rect 9928 4868 9932 4924
rect 9932 4868 9988 4924
rect 9988 4868 9992 4924
rect 9928 4864 9992 4868
rect 10008 4924 10072 4928
rect 10008 4868 10012 4924
rect 10012 4868 10068 4924
rect 10068 4868 10072 4924
rect 10008 4864 10072 4868
rect 10088 4924 10152 4928
rect 10088 4868 10092 4924
rect 10092 4868 10148 4924
rect 10148 4868 10152 4924
rect 10088 4864 10152 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 15938 4924 16002 4928
rect 15938 4868 15942 4924
rect 15942 4868 15998 4924
rect 15998 4868 16002 4924
rect 15938 4864 16002 4868
rect 16018 4924 16082 4928
rect 16018 4868 16022 4924
rect 16022 4868 16078 4924
rect 16078 4868 16082 4924
rect 16018 4864 16082 4868
rect 6882 4380 6946 4384
rect 6882 4324 6886 4380
rect 6886 4324 6942 4380
rect 6942 4324 6946 4380
rect 6882 4320 6946 4324
rect 6962 4380 7026 4384
rect 6962 4324 6966 4380
rect 6966 4324 7022 4380
rect 7022 4324 7026 4380
rect 6962 4320 7026 4324
rect 7042 4380 7106 4384
rect 7042 4324 7046 4380
rect 7046 4324 7102 4380
rect 7102 4324 7106 4380
rect 7042 4320 7106 4324
rect 7122 4380 7186 4384
rect 7122 4324 7126 4380
rect 7126 4324 7182 4380
rect 7182 4324 7186 4380
rect 7122 4320 7186 4324
rect 12813 4380 12877 4384
rect 12813 4324 12817 4380
rect 12817 4324 12873 4380
rect 12873 4324 12877 4380
rect 12813 4320 12877 4324
rect 12893 4380 12957 4384
rect 12893 4324 12897 4380
rect 12897 4324 12953 4380
rect 12953 4324 12957 4380
rect 12893 4320 12957 4324
rect 12973 4380 13037 4384
rect 12973 4324 12977 4380
rect 12977 4324 13033 4380
rect 13033 4324 13037 4380
rect 12973 4320 13037 4324
rect 13053 4380 13117 4384
rect 13053 4324 13057 4380
rect 13057 4324 13113 4380
rect 13113 4324 13117 4380
rect 13053 4320 13117 4324
rect 3917 3836 3981 3840
rect 3917 3780 3921 3836
rect 3921 3780 3977 3836
rect 3977 3780 3981 3836
rect 3917 3776 3981 3780
rect 3997 3836 4061 3840
rect 3997 3780 4001 3836
rect 4001 3780 4057 3836
rect 4057 3780 4061 3836
rect 3997 3776 4061 3780
rect 4077 3836 4141 3840
rect 4077 3780 4081 3836
rect 4081 3780 4137 3836
rect 4137 3780 4141 3836
rect 4077 3776 4141 3780
rect 4157 3836 4221 3840
rect 4157 3780 4161 3836
rect 4161 3780 4217 3836
rect 4217 3780 4221 3836
rect 4157 3776 4221 3780
rect 9848 3836 9912 3840
rect 9848 3780 9852 3836
rect 9852 3780 9908 3836
rect 9908 3780 9912 3836
rect 9848 3776 9912 3780
rect 9928 3836 9992 3840
rect 9928 3780 9932 3836
rect 9932 3780 9988 3836
rect 9988 3780 9992 3836
rect 9928 3776 9992 3780
rect 10008 3836 10072 3840
rect 10008 3780 10012 3836
rect 10012 3780 10068 3836
rect 10068 3780 10072 3836
rect 10008 3776 10072 3780
rect 10088 3836 10152 3840
rect 10088 3780 10092 3836
rect 10092 3780 10148 3836
rect 10148 3780 10152 3836
rect 10088 3776 10152 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 15938 3836 16002 3840
rect 15938 3780 15942 3836
rect 15942 3780 15998 3836
rect 15998 3780 16002 3836
rect 15938 3776 16002 3780
rect 16018 3836 16082 3840
rect 16018 3780 16022 3836
rect 16022 3780 16078 3836
rect 16078 3780 16082 3836
rect 16018 3776 16082 3780
rect 6882 3292 6946 3296
rect 6882 3236 6886 3292
rect 6886 3236 6942 3292
rect 6942 3236 6946 3292
rect 6882 3232 6946 3236
rect 6962 3292 7026 3296
rect 6962 3236 6966 3292
rect 6966 3236 7022 3292
rect 7022 3236 7026 3292
rect 6962 3232 7026 3236
rect 7042 3292 7106 3296
rect 7042 3236 7046 3292
rect 7046 3236 7102 3292
rect 7102 3236 7106 3292
rect 7042 3232 7106 3236
rect 7122 3292 7186 3296
rect 7122 3236 7126 3292
rect 7126 3236 7182 3292
rect 7182 3236 7186 3292
rect 7122 3232 7186 3236
rect 12813 3292 12877 3296
rect 12813 3236 12817 3292
rect 12817 3236 12873 3292
rect 12873 3236 12877 3292
rect 12813 3232 12877 3236
rect 12893 3292 12957 3296
rect 12893 3236 12897 3292
rect 12897 3236 12953 3292
rect 12953 3236 12957 3292
rect 12893 3232 12957 3236
rect 12973 3292 13037 3296
rect 12973 3236 12977 3292
rect 12977 3236 13033 3292
rect 13033 3236 13037 3292
rect 12973 3232 13037 3236
rect 13053 3292 13117 3296
rect 13053 3236 13057 3292
rect 13057 3236 13113 3292
rect 13113 3236 13117 3292
rect 13053 3232 13117 3236
rect 3917 2748 3981 2752
rect 3917 2692 3921 2748
rect 3921 2692 3977 2748
rect 3977 2692 3981 2748
rect 3917 2688 3981 2692
rect 3997 2748 4061 2752
rect 3997 2692 4001 2748
rect 4001 2692 4057 2748
rect 4057 2692 4061 2748
rect 3997 2688 4061 2692
rect 4077 2748 4141 2752
rect 4077 2692 4081 2748
rect 4081 2692 4137 2748
rect 4137 2692 4141 2748
rect 4077 2688 4141 2692
rect 4157 2748 4221 2752
rect 4157 2692 4161 2748
rect 4161 2692 4217 2748
rect 4217 2692 4221 2748
rect 4157 2688 4221 2692
rect 9848 2748 9912 2752
rect 9848 2692 9852 2748
rect 9852 2692 9908 2748
rect 9908 2692 9912 2748
rect 9848 2688 9912 2692
rect 9928 2748 9992 2752
rect 9928 2692 9932 2748
rect 9932 2692 9988 2748
rect 9988 2692 9992 2748
rect 9928 2688 9992 2692
rect 10008 2748 10072 2752
rect 10008 2692 10012 2748
rect 10012 2692 10068 2748
rect 10068 2692 10072 2748
rect 10008 2688 10072 2692
rect 10088 2748 10152 2752
rect 10088 2692 10092 2748
rect 10092 2692 10148 2748
rect 10148 2692 10152 2748
rect 10088 2688 10152 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 15938 2748 16002 2752
rect 15938 2692 15942 2748
rect 15942 2692 15998 2748
rect 15998 2692 16002 2748
rect 15938 2688 16002 2692
rect 16018 2748 16082 2752
rect 16018 2692 16022 2748
rect 16022 2692 16078 2748
rect 16078 2692 16082 2748
rect 16018 2688 16082 2692
rect 6882 2204 6946 2208
rect 6882 2148 6886 2204
rect 6886 2148 6942 2204
rect 6942 2148 6946 2204
rect 6882 2144 6946 2148
rect 6962 2204 7026 2208
rect 6962 2148 6966 2204
rect 6966 2148 7022 2204
rect 7022 2148 7026 2204
rect 6962 2144 7026 2148
rect 7042 2204 7106 2208
rect 7042 2148 7046 2204
rect 7046 2148 7102 2204
rect 7102 2148 7106 2204
rect 7042 2144 7106 2148
rect 7122 2204 7186 2208
rect 7122 2148 7126 2204
rect 7126 2148 7182 2204
rect 7182 2148 7186 2204
rect 7122 2144 7186 2148
rect 12813 2204 12877 2208
rect 12813 2148 12817 2204
rect 12817 2148 12873 2204
rect 12873 2148 12877 2204
rect 12813 2144 12877 2148
rect 12893 2204 12957 2208
rect 12893 2148 12897 2204
rect 12897 2148 12953 2204
rect 12953 2148 12957 2204
rect 12893 2144 12957 2148
rect 12973 2204 13037 2208
rect 12973 2148 12977 2204
rect 12977 2148 13033 2204
rect 13033 2148 13037 2204
rect 12973 2144 13037 2148
rect 13053 2204 13117 2208
rect 13053 2148 13057 2204
rect 13057 2148 13113 2204
rect 13113 2148 13117 2204
rect 13053 2144 13117 2148
<< metal4 >>
rect 3909 47360 4230 47376
rect 3909 47296 3917 47360
rect 3981 47296 3997 47360
rect 4061 47296 4077 47360
rect 4141 47296 4157 47360
rect 4221 47296 4230 47360
rect 3909 46272 4230 47296
rect 3909 46208 3917 46272
rect 3981 46208 3997 46272
rect 4061 46208 4077 46272
rect 4141 46208 4157 46272
rect 4221 46208 4230 46272
rect 3909 45184 4230 46208
rect 3909 45120 3917 45184
rect 3981 45120 3997 45184
rect 4061 45120 4077 45184
rect 4141 45120 4157 45184
rect 4221 45120 4230 45184
rect 3909 44096 4230 45120
rect 3909 44032 3917 44096
rect 3981 44032 3997 44096
rect 4061 44032 4077 44096
rect 4141 44032 4157 44096
rect 4221 44032 4230 44096
rect 3909 43008 4230 44032
rect 3909 42944 3917 43008
rect 3981 42944 3997 43008
rect 4061 42944 4077 43008
rect 4141 42944 4157 43008
rect 4221 42944 4230 43008
rect 3909 41920 4230 42944
rect 3909 41856 3917 41920
rect 3981 41856 3997 41920
rect 4061 41856 4077 41920
rect 4141 41856 4157 41920
rect 4221 41856 4230 41920
rect 3909 40832 4230 41856
rect 3909 40768 3917 40832
rect 3981 40768 3997 40832
rect 4061 40768 4077 40832
rect 4141 40768 4157 40832
rect 4221 40768 4230 40832
rect 3909 39744 4230 40768
rect 3909 39680 3917 39744
rect 3981 39680 3997 39744
rect 4061 39680 4077 39744
rect 4141 39680 4157 39744
rect 4221 39680 4230 39744
rect 3909 38656 4230 39680
rect 3909 38592 3917 38656
rect 3981 38592 3997 38656
rect 4061 38592 4077 38656
rect 4141 38592 4157 38656
rect 4221 38592 4230 38656
rect 3909 37568 4230 38592
rect 3909 37504 3917 37568
rect 3981 37504 3997 37568
rect 4061 37504 4077 37568
rect 4141 37504 4157 37568
rect 4221 37504 4230 37568
rect 3909 36480 4230 37504
rect 3909 36416 3917 36480
rect 3981 36416 3997 36480
rect 4061 36416 4077 36480
rect 4141 36416 4157 36480
rect 4221 36416 4230 36480
rect 3909 35392 4230 36416
rect 3909 35328 3917 35392
rect 3981 35328 3997 35392
rect 4061 35328 4077 35392
rect 4141 35328 4157 35392
rect 4221 35328 4230 35392
rect 3909 34304 4230 35328
rect 3909 34240 3917 34304
rect 3981 34240 3997 34304
rect 4061 34240 4077 34304
rect 4141 34240 4157 34304
rect 4221 34240 4230 34304
rect 3909 33216 4230 34240
rect 3909 33152 3917 33216
rect 3981 33152 3997 33216
rect 4061 33152 4077 33216
rect 4141 33152 4157 33216
rect 4221 33152 4230 33216
rect 3909 32128 4230 33152
rect 3909 32064 3917 32128
rect 3981 32064 3997 32128
rect 4061 32064 4077 32128
rect 4141 32064 4157 32128
rect 4221 32064 4230 32128
rect 3909 31040 4230 32064
rect 3909 30976 3917 31040
rect 3981 30976 3997 31040
rect 4061 30976 4077 31040
rect 4141 30976 4157 31040
rect 4221 30976 4230 31040
rect 3909 29952 4230 30976
rect 3909 29888 3917 29952
rect 3981 29888 3997 29952
rect 4061 29888 4077 29952
rect 4141 29888 4157 29952
rect 4221 29888 4230 29952
rect 3909 28864 4230 29888
rect 3909 28800 3917 28864
rect 3981 28800 3997 28864
rect 4061 28800 4077 28864
rect 4141 28800 4157 28864
rect 4221 28800 4230 28864
rect 3909 27776 4230 28800
rect 3909 27712 3917 27776
rect 3981 27712 3997 27776
rect 4061 27712 4077 27776
rect 4141 27712 4157 27776
rect 4221 27712 4230 27776
rect 3909 26688 4230 27712
rect 3909 26624 3917 26688
rect 3981 26624 3997 26688
rect 4061 26624 4077 26688
rect 4141 26624 4157 26688
rect 4221 26624 4230 26688
rect 3909 25600 4230 26624
rect 3909 25536 3917 25600
rect 3981 25536 3997 25600
rect 4061 25536 4077 25600
rect 4141 25536 4157 25600
rect 4221 25536 4230 25600
rect 3909 24512 4230 25536
rect 3909 24448 3917 24512
rect 3981 24448 3997 24512
rect 4061 24448 4077 24512
rect 4141 24448 4157 24512
rect 4221 24448 4230 24512
rect 3909 23424 4230 24448
rect 3909 23360 3917 23424
rect 3981 23360 3997 23424
rect 4061 23360 4077 23424
rect 4141 23360 4157 23424
rect 4221 23360 4230 23424
rect 3909 22336 4230 23360
rect 3909 22272 3917 22336
rect 3981 22272 3997 22336
rect 4061 22272 4077 22336
rect 4141 22272 4157 22336
rect 4221 22272 4230 22336
rect 3909 21248 4230 22272
rect 3909 21184 3917 21248
rect 3981 21184 3997 21248
rect 4061 21184 4077 21248
rect 4141 21184 4157 21248
rect 4221 21184 4230 21248
rect 3909 20160 4230 21184
rect 3909 20096 3917 20160
rect 3981 20096 3997 20160
rect 4061 20096 4077 20160
rect 4141 20096 4157 20160
rect 4221 20096 4230 20160
rect 3909 19072 4230 20096
rect 3909 19008 3917 19072
rect 3981 19008 3997 19072
rect 4061 19008 4077 19072
rect 4141 19008 4157 19072
rect 4221 19008 4230 19072
rect 3909 17984 4230 19008
rect 3909 17920 3917 17984
rect 3981 17920 3997 17984
rect 4061 17920 4077 17984
rect 4141 17920 4157 17984
rect 4221 17920 4230 17984
rect 3909 16896 4230 17920
rect 3909 16832 3917 16896
rect 3981 16832 3997 16896
rect 4061 16832 4077 16896
rect 4141 16832 4157 16896
rect 4221 16832 4230 16896
rect 3909 15808 4230 16832
rect 3909 15744 3917 15808
rect 3981 15744 3997 15808
rect 4061 15744 4077 15808
rect 4141 15744 4157 15808
rect 4221 15744 4230 15808
rect 3909 14720 4230 15744
rect 3909 14656 3917 14720
rect 3981 14656 3997 14720
rect 4061 14656 4077 14720
rect 4141 14656 4157 14720
rect 4221 14656 4230 14720
rect 3909 13632 4230 14656
rect 3909 13568 3917 13632
rect 3981 13568 3997 13632
rect 4061 13568 4077 13632
rect 4141 13568 4157 13632
rect 4221 13568 4230 13632
rect 3909 12544 4230 13568
rect 3909 12480 3917 12544
rect 3981 12480 3997 12544
rect 4061 12480 4077 12544
rect 4141 12480 4157 12544
rect 4221 12480 4230 12544
rect 3909 11456 4230 12480
rect 3909 11392 3917 11456
rect 3981 11392 3997 11456
rect 4061 11392 4077 11456
rect 4141 11392 4157 11456
rect 4221 11392 4230 11456
rect 3909 10368 4230 11392
rect 3909 10304 3917 10368
rect 3981 10304 3997 10368
rect 4061 10304 4077 10368
rect 4141 10304 4157 10368
rect 4221 10304 4230 10368
rect 3909 9280 4230 10304
rect 3909 9216 3917 9280
rect 3981 9216 3997 9280
rect 4061 9216 4077 9280
rect 4141 9216 4157 9280
rect 4221 9216 4230 9280
rect 3909 8192 4230 9216
rect 3909 8128 3917 8192
rect 3981 8128 3997 8192
rect 4061 8128 4077 8192
rect 4141 8128 4157 8192
rect 4221 8128 4230 8192
rect 3909 7104 4230 8128
rect 3909 7040 3917 7104
rect 3981 7040 3997 7104
rect 4061 7040 4077 7104
rect 4141 7040 4157 7104
rect 4221 7040 4230 7104
rect 3909 6016 4230 7040
rect 3909 5952 3917 6016
rect 3981 5952 3997 6016
rect 4061 5952 4077 6016
rect 4141 5952 4157 6016
rect 4221 5952 4230 6016
rect 3909 4928 4230 5952
rect 3909 4864 3917 4928
rect 3981 4864 3997 4928
rect 4061 4864 4077 4928
rect 4141 4864 4157 4928
rect 4221 4864 4230 4928
rect 3909 3840 4230 4864
rect 3909 3776 3917 3840
rect 3981 3776 3997 3840
rect 4061 3776 4077 3840
rect 4141 3776 4157 3840
rect 4221 3776 4230 3840
rect 3909 2752 4230 3776
rect 3909 2688 3917 2752
rect 3981 2688 3997 2752
rect 4061 2688 4077 2752
rect 4141 2688 4157 2752
rect 4221 2688 4230 2752
rect 3909 2128 4230 2688
rect 6874 46816 7194 47376
rect 6874 46752 6882 46816
rect 6946 46752 6962 46816
rect 7026 46752 7042 46816
rect 7106 46752 7122 46816
rect 7186 46752 7194 46816
rect 6874 45728 7194 46752
rect 6874 45664 6882 45728
rect 6946 45664 6962 45728
rect 7026 45664 7042 45728
rect 7106 45664 7122 45728
rect 7186 45664 7194 45728
rect 6874 44640 7194 45664
rect 6874 44576 6882 44640
rect 6946 44576 6962 44640
rect 7026 44576 7042 44640
rect 7106 44576 7122 44640
rect 7186 44576 7194 44640
rect 6874 43552 7194 44576
rect 6874 43488 6882 43552
rect 6946 43488 6962 43552
rect 7026 43488 7042 43552
rect 7106 43488 7122 43552
rect 7186 43488 7194 43552
rect 6874 42464 7194 43488
rect 6874 42400 6882 42464
rect 6946 42400 6962 42464
rect 7026 42400 7042 42464
rect 7106 42400 7122 42464
rect 7186 42400 7194 42464
rect 6874 41376 7194 42400
rect 6874 41312 6882 41376
rect 6946 41312 6962 41376
rect 7026 41312 7042 41376
rect 7106 41312 7122 41376
rect 7186 41312 7194 41376
rect 6874 40288 7194 41312
rect 6874 40224 6882 40288
rect 6946 40224 6962 40288
rect 7026 40224 7042 40288
rect 7106 40224 7122 40288
rect 7186 40224 7194 40288
rect 6874 39200 7194 40224
rect 6874 39136 6882 39200
rect 6946 39136 6962 39200
rect 7026 39136 7042 39200
rect 7106 39136 7122 39200
rect 7186 39136 7194 39200
rect 6874 38112 7194 39136
rect 6874 38048 6882 38112
rect 6946 38048 6962 38112
rect 7026 38048 7042 38112
rect 7106 38048 7122 38112
rect 7186 38048 7194 38112
rect 6874 37024 7194 38048
rect 6874 36960 6882 37024
rect 6946 36960 6962 37024
rect 7026 36960 7042 37024
rect 7106 36960 7122 37024
rect 7186 36960 7194 37024
rect 6874 35936 7194 36960
rect 6874 35872 6882 35936
rect 6946 35872 6962 35936
rect 7026 35872 7042 35936
rect 7106 35872 7122 35936
rect 7186 35872 7194 35936
rect 6874 34848 7194 35872
rect 6874 34784 6882 34848
rect 6946 34784 6962 34848
rect 7026 34784 7042 34848
rect 7106 34784 7122 34848
rect 7186 34784 7194 34848
rect 6874 33760 7194 34784
rect 6874 33696 6882 33760
rect 6946 33696 6962 33760
rect 7026 33696 7042 33760
rect 7106 33696 7122 33760
rect 7186 33696 7194 33760
rect 6874 32672 7194 33696
rect 6874 32608 6882 32672
rect 6946 32608 6962 32672
rect 7026 32608 7042 32672
rect 7106 32608 7122 32672
rect 7186 32608 7194 32672
rect 6874 31584 7194 32608
rect 6874 31520 6882 31584
rect 6946 31520 6962 31584
rect 7026 31520 7042 31584
rect 7106 31520 7122 31584
rect 7186 31520 7194 31584
rect 6874 30496 7194 31520
rect 6874 30432 6882 30496
rect 6946 30432 6962 30496
rect 7026 30432 7042 30496
rect 7106 30432 7122 30496
rect 7186 30432 7194 30496
rect 6874 29408 7194 30432
rect 6874 29344 6882 29408
rect 6946 29344 6962 29408
rect 7026 29344 7042 29408
rect 7106 29344 7122 29408
rect 7186 29344 7194 29408
rect 6874 28320 7194 29344
rect 6874 28256 6882 28320
rect 6946 28256 6962 28320
rect 7026 28256 7042 28320
rect 7106 28256 7122 28320
rect 7186 28256 7194 28320
rect 6874 27232 7194 28256
rect 6874 27168 6882 27232
rect 6946 27168 6962 27232
rect 7026 27168 7042 27232
rect 7106 27168 7122 27232
rect 7186 27168 7194 27232
rect 6874 26144 7194 27168
rect 6874 26080 6882 26144
rect 6946 26080 6962 26144
rect 7026 26080 7042 26144
rect 7106 26080 7122 26144
rect 7186 26080 7194 26144
rect 6874 25056 7194 26080
rect 6874 24992 6882 25056
rect 6946 24992 6962 25056
rect 7026 24992 7042 25056
rect 7106 24992 7122 25056
rect 7186 24992 7194 25056
rect 6874 23968 7194 24992
rect 6874 23904 6882 23968
rect 6946 23904 6962 23968
rect 7026 23904 7042 23968
rect 7106 23904 7122 23968
rect 7186 23904 7194 23968
rect 6874 22880 7194 23904
rect 6874 22816 6882 22880
rect 6946 22816 6962 22880
rect 7026 22816 7042 22880
rect 7106 22816 7122 22880
rect 7186 22816 7194 22880
rect 6874 21792 7194 22816
rect 6874 21728 6882 21792
rect 6946 21728 6962 21792
rect 7026 21728 7042 21792
rect 7106 21728 7122 21792
rect 7186 21728 7194 21792
rect 6874 20704 7194 21728
rect 6874 20640 6882 20704
rect 6946 20640 6962 20704
rect 7026 20640 7042 20704
rect 7106 20640 7122 20704
rect 7186 20640 7194 20704
rect 6874 19616 7194 20640
rect 6874 19552 6882 19616
rect 6946 19552 6962 19616
rect 7026 19552 7042 19616
rect 7106 19552 7122 19616
rect 7186 19552 7194 19616
rect 6874 18528 7194 19552
rect 6874 18464 6882 18528
rect 6946 18464 6962 18528
rect 7026 18464 7042 18528
rect 7106 18464 7122 18528
rect 7186 18464 7194 18528
rect 6874 17440 7194 18464
rect 6874 17376 6882 17440
rect 6946 17376 6962 17440
rect 7026 17376 7042 17440
rect 7106 17376 7122 17440
rect 7186 17376 7194 17440
rect 6874 16352 7194 17376
rect 6874 16288 6882 16352
rect 6946 16288 6962 16352
rect 7026 16288 7042 16352
rect 7106 16288 7122 16352
rect 7186 16288 7194 16352
rect 6874 15264 7194 16288
rect 6874 15200 6882 15264
rect 6946 15200 6962 15264
rect 7026 15200 7042 15264
rect 7106 15200 7122 15264
rect 7186 15200 7194 15264
rect 6874 14176 7194 15200
rect 6874 14112 6882 14176
rect 6946 14112 6962 14176
rect 7026 14112 7042 14176
rect 7106 14112 7122 14176
rect 7186 14112 7194 14176
rect 6874 13088 7194 14112
rect 6874 13024 6882 13088
rect 6946 13024 6962 13088
rect 7026 13024 7042 13088
rect 7106 13024 7122 13088
rect 7186 13024 7194 13088
rect 6874 12000 7194 13024
rect 6874 11936 6882 12000
rect 6946 11936 6962 12000
rect 7026 11936 7042 12000
rect 7106 11936 7122 12000
rect 7186 11936 7194 12000
rect 6874 10912 7194 11936
rect 6874 10848 6882 10912
rect 6946 10848 6962 10912
rect 7026 10848 7042 10912
rect 7106 10848 7122 10912
rect 7186 10848 7194 10912
rect 6874 9824 7194 10848
rect 6874 9760 6882 9824
rect 6946 9760 6962 9824
rect 7026 9760 7042 9824
rect 7106 9760 7122 9824
rect 7186 9760 7194 9824
rect 6874 8736 7194 9760
rect 6874 8672 6882 8736
rect 6946 8672 6962 8736
rect 7026 8672 7042 8736
rect 7106 8672 7122 8736
rect 7186 8672 7194 8736
rect 6874 7648 7194 8672
rect 6874 7584 6882 7648
rect 6946 7584 6962 7648
rect 7026 7584 7042 7648
rect 7106 7584 7122 7648
rect 7186 7584 7194 7648
rect 6874 6560 7194 7584
rect 6874 6496 6882 6560
rect 6946 6496 6962 6560
rect 7026 6496 7042 6560
rect 7106 6496 7122 6560
rect 7186 6496 7194 6560
rect 6874 5472 7194 6496
rect 6874 5408 6882 5472
rect 6946 5408 6962 5472
rect 7026 5408 7042 5472
rect 7106 5408 7122 5472
rect 7186 5408 7194 5472
rect 6874 4384 7194 5408
rect 6874 4320 6882 4384
rect 6946 4320 6962 4384
rect 7026 4320 7042 4384
rect 7106 4320 7122 4384
rect 7186 4320 7194 4384
rect 6874 3296 7194 4320
rect 6874 3232 6882 3296
rect 6946 3232 6962 3296
rect 7026 3232 7042 3296
rect 7106 3232 7122 3296
rect 7186 3232 7194 3296
rect 6874 2208 7194 3232
rect 6874 2144 6882 2208
rect 6946 2144 6962 2208
rect 7026 2144 7042 2208
rect 7106 2144 7122 2208
rect 7186 2144 7194 2208
rect 6874 2128 7194 2144
rect 9840 47360 10160 47376
rect 9840 47296 9848 47360
rect 9912 47296 9928 47360
rect 9992 47296 10008 47360
rect 10072 47296 10088 47360
rect 10152 47296 10160 47360
rect 9840 46272 10160 47296
rect 9840 46208 9848 46272
rect 9912 46208 9928 46272
rect 9992 46208 10008 46272
rect 10072 46208 10088 46272
rect 10152 46208 10160 46272
rect 9840 45184 10160 46208
rect 9840 45120 9848 45184
rect 9912 45120 9928 45184
rect 9992 45120 10008 45184
rect 10072 45120 10088 45184
rect 10152 45120 10160 45184
rect 9840 44096 10160 45120
rect 9840 44032 9848 44096
rect 9912 44032 9928 44096
rect 9992 44032 10008 44096
rect 10072 44032 10088 44096
rect 10152 44032 10160 44096
rect 9840 43008 10160 44032
rect 9840 42944 9848 43008
rect 9912 42944 9928 43008
rect 9992 42944 10008 43008
rect 10072 42944 10088 43008
rect 10152 42944 10160 43008
rect 9840 41920 10160 42944
rect 9840 41856 9848 41920
rect 9912 41856 9928 41920
rect 9992 41856 10008 41920
rect 10072 41856 10088 41920
rect 10152 41856 10160 41920
rect 9840 40832 10160 41856
rect 9840 40768 9848 40832
rect 9912 40768 9928 40832
rect 9992 40768 10008 40832
rect 10072 40768 10088 40832
rect 10152 40768 10160 40832
rect 9840 39744 10160 40768
rect 9840 39680 9848 39744
rect 9912 39680 9928 39744
rect 9992 39680 10008 39744
rect 10072 39680 10088 39744
rect 10152 39680 10160 39744
rect 9840 38656 10160 39680
rect 9840 38592 9848 38656
rect 9912 38592 9928 38656
rect 9992 38592 10008 38656
rect 10072 38592 10088 38656
rect 10152 38592 10160 38656
rect 9840 37568 10160 38592
rect 9840 37504 9848 37568
rect 9912 37504 9928 37568
rect 9992 37504 10008 37568
rect 10072 37504 10088 37568
rect 10152 37504 10160 37568
rect 9840 36480 10160 37504
rect 9840 36416 9848 36480
rect 9912 36416 9928 36480
rect 9992 36416 10008 36480
rect 10072 36416 10088 36480
rect 10152 36416 10160 36480
rect 9840 35392 10160 36416
rect 9840 35328 9848 35392
rect 9912 35328 9928 35392
rect 9992 35328 10008 35392
rect 10072 35328 10088 35392
rect 10152 35328 10160 35392
rect 9840 34304 10160 35328
rect 9840 34240 9848 34304
rect 9912 34240 9928 34304
rect 9992 34240 10008 34304
rect 10072 34240 10088 34304
rect 10152 34240 10160 34304
rect 9840 33216 10160 34240
rect 9840 33152 9848 33216
rect 9912 33152 9928 33216
rect 9992 33152 10008 33216
rect 10072 33152 10088 33216
rect 10152 33152 10160 33216
rect 9840 32128 10160 33152
rect 9840 32064 9848 32128
rect 9912 32064 9928 32128
rect 9992 32064 10008 32128
rect 10072 32064 10088 32128
rect 10152 32064 10160 32128
rect 9840 31040 10160 32064
rect 9840 30976 9848 31040
rect 9912 30976 9928 31040
rect 9992 30976 10008 31040
rect 10072 30976 10088 31040
rect 10152 30976 10160 31040
rect 9840 29952 10160 30976
rect 9840 29888 9848 29952
rect 9912 29888 9928 29952
rect 9992 29888 10008 29952
rect 10072 29888 10088 29952
rect 10152 29888 10160 29952
rect 9840 28864 10160 29888
rect 9840 28800 9848 28864
rect 9912 28800 9928 28864
rect 9992 28800 10008 28864
rect 10072 28800 10088 28864
rect 10152 28800 10160 28864
rect 9840 27776 10160 28800
rect 9840 27712 9848 27776
rect 9912 27712 9928 27776
rect 9992 27712 10008 27776
rect 10072 27712 10088 27776
rect 10152 27712 10160 27776
rect 9840 26688 10160 27712
rect 9840 26624 9848 26688
rect 9912 26624 9928 26688
rect 9992 26624 10008 26688
rect 10072 26624 10088 26688
rect 10152 26624 10160 26688
rect 9840 25600 10160 26624
rect 9840 25536 9848 25600
rect 9912 25536 9928 25600
rect 9992 25536 10008 25600
rect 10072 25536 10088 25600
rect 10152 25536 10160 25600
rect 9840 24512 10160 25536
rect 9840 24448 9848 24512
rect 9912 24448 9928 24512
rect 9992 24448 10008 24512
rect 10072 24448 10088 24512
rect 10152 24448 10160 24512
rect 9840 23424 10160 24448
rect 9840 23360 9848 23424
rect 9912 23360 9928 23424
rect 9992 23360 10008 23424
rect 10072 23360 10088 23424
rect 10152 23360 10160 23424
rect 9840 22336 10160 23360
rect 9840 22272 9848 22336
rect 9912 22272 9928 22336
rect 9992 22272 10008 22336
rect 10072 22272 10088 22336
rect 10152 22272 10160 22336
rect 9840 21248 10160 22272
rect 9840 21184 9848 21248
rect 9912 21184 9928 21248
rect 9992 21184 10008 21248
rect 10072 21184 10088 21248
rect 10152 21184 10160 21248
rect 9840 20160 10160 21184
rect 9840 20096 9848 20160
rect 9912 20096 9928 20160
rect 9992 20096 10008 20160
rect 10072 20096 10088 20160
rect 10152 20096 10160 20160
rect 9840 19072 10160 20096
rect 9840 19008 9848 19072
rect 9912 19008 9928 19072
rect 9992 19008 10008 19072
rect 10072 19008 10088 19072
rect 10152 19008 10160 19072
rect 9840 17984 10160 19008
rect 9840 17920 9848 17984
rect 9912 17920 9928 17984
rect 9992 17920 10008 17984
rect 10072 17920 10088 17984
rect 10152 17920 10160 17984
rect 9840 16896 10160 17920
rect 9840 16832 9848 16896
rect 9912 16832 9928 16896
rect 9992 16832 10008 16896
rect 10072 16832 10088 16896
rect 10152 16832 10160 16896
rect 9840 15808 10160 16832
rect 9840 15744 9848 15808
rect 9912 15744 9928 15808
rect 9992 15744 10008 15808
rect 10072 15744 10088 15808
rect 10152 15744 10160 15808
rect 9840 14720 10160 15744
rect 9840 14656 9848 14720
rect 9912 14656 9928 14720
rect 9992 14656 10008 14720
rect 10072 14656 10088 14720
rect 10152 14656 10160 14720
rect 9840 13632 10160 14656
rect 9840 13568 9848 13632
rect 9912 13568 9928 13632
rect 9992 13568 10008 13632
rect 10072 13568 10088 13632
rect 10152 13568 10160 13632
rect 9840 12544 10160 13568
rect 9840 12480 9848 12544
rect 9912 12480 9928 12544
rect 9992 12480 10008 12544
rect 10072 12480 10088 12544
rect 10152 12480 10160 12544
rect 9840 11456 10160 12480
rect 9840 11392 9848 11456
rect 9912 11392 9928 11456
rect 9992 11392 10008 11456
rect 10072 11392 10088 11456
rect 10152 11392 10160 11456
rect 9840 10368 10160 11392
rect 9840 10304 9848 10368
rect 9912 10304 9928 10368
rect 9992 10304 10008 10368
rect 10072 10304 10088 10368
rect 10152 10304 10160 10368
rect 9840 9280 10160 10304
rect 9840 9216 9848 9280
rect 9912 9216 9928 9280
rect 9992 9216 10008 9280
rect 10072 9216 10088 9280
rect 10152 9216 10160 9280
rect 9840 8192 10160 9216
rect 9840 8128 9848 8192
rect 9912 8128 9928 8192
rect 9992 8128 10008 8192
rect 10072 8128 10088 8192
rect 10152 8128 10160 8192
rect 9840 7104 10160 8128
rect 9840 7040 9848 7104
rect 9912 7040 9928 7104
rect 9992 7040 10008 7104
rect 10072 7040 10088 7104
rect 10152 7040 10160 7104
rect 9840 6016 10160 7040
rect 9840 5952 9848 6016
rect 9912 5952 9928 6016
rect 9992 5952 10008 6016
rect 10072 5952 10088 6016
rect 10152 5952 10160 6016
rect 9840 4928 10160 5952
rect 9840 4864 9848 4928
rect 9912 4864 9928 4928
rect 9992 4864 10008 4928
rect 10072 4864 10088 4928
rect 10152 4864 10160 4928
rect 9840 3840 10160 4864
rect 9840 3776 9848 3840
rect 9912 3776 9928 3840
rect 9992 3776 10008 3840
rect 10072 3776 10088 3840
rect 10152 3776 10160 3840
rect 9840 2752 10160 3776
rect 9840 2688 9848 2752
rect 9912 2688 9928 2752
rect 9992 2688 10008 2752
rect 10072 2688 10088 2752
rect 10152 2688 10160 2752
rect 9840 2128 10160 2688
rect 12805 46816 13125 47376
rect 12805 46752 12813 46816
rect 12877 46752 12893 46816
rect 12957 46752 12973 46816
rect 13037 46752 13053 46816
rect 13117 46752 13125 46816
rect 12805 45728 13125 46752
rect 12805 45664 12813 45728
rect 12877 45664 12893 45728
rect 12957 45664 12973 45728
rect 13037 45664 13053 45728
rect 13117 45664 13125 45728
rect 12805 44640 13125 45664
rect 12805 44576 12813 44640
rect 12877 44576 12893 44640
rect 12957 44576 12973 44640
rect 13037 44576 13053 44640
rect 13117 44576 13125 44640
rect 12805 43552 13125 44576
rect 12805 43488 12813 43552
rect 12877 43488 12893 43552
rect 12957 43488 12973 43552
rect 13037 43488 13053 43552
rect 13117 43488 13125 43552
rect 12805 42464 13125 43488
rect 12805 42400 12813 42464
rect 12877 42400 12893 42464
rect 12957 42400 12973 42464
rect 13037 42400 13053 42464
rect 13117 42400 13125 42464
rect 12805 41376 13125 42400
rect 12805 41312 12813 41376
rect 12877 41312 12893 41376
rect 12957 41312 12973 41376
rect 13037 41312 13053 41376
rect 13117 41312 13125 41376
rect 12805 40288 13125 41312
rect 12805 40224 12813 40288
rect 12877 40224 12893 40288
rect 12957 40224 12973 40288
rect 13037 40224 13053 40288
rect 13117 40224 13125 40288
rect 12805 39200 13125 40224
rect 12805 39136 12813 39200
rect 12877 39136 12893 39200
rect 12957 39136 12973 39200
rect 13037 39136 13053 39200
rect 13117 39136 13125 39200
rect 12805 38112 13125 39136
rect 12805 38048 12813 38112
rect 12877 38048 12893 38112
rect 12957 38048 12973 38112
rect 13037 38048 13053 38112
rect 13117 38048 13125 38112
rect 12805 37024 13125 38048
rect 12805 36960 12813 37024
rect 12877 36960 12893 37024
rect 12957 36960 12973 37024
rect 13037 36960 13053 37024
rect 13117 36960 13125 37024
rect 12805 35936 13125 36960
rect 12805 35872 12813 35936
rect 12877 35872 12893 35936
rect 12957 35872 12973 35936
rect 13037 35872 13053 35936
rect 13117 35872 13125 35936
rect 12805 34848 13125 35872
rect 12805 34784 12813 34848
rect 12877 34784 12893 34848
rect 12957 34784 12973 34848
rect 13037 34784 13053 34848
rect 13117 34784 13125 34848
rect 12805 33760 13125 34784
rect 12805 33696 12813 33760
rect 12877 33696 12893 33760
rect 12957 33696 12973 33760
rect 13037 33696 13053 33760
rect 13117 33696 13125 33760
rect 12805 32672 13125 33696
rect 12805 32608 12813 32672
rect 12877 32608 12893 32672
rect 12957 32608 12973 32672
rect 13037 32608 13053 32672
rect 13117 32608 13125 32672
rect 12805 31584 13125 32608
rect 12805 31520 12813 31584
rect 12877 31520 12893 31584
rect 12957 31520 12973 31584
rect 13037 31520 13053 31584
rect 13117 31520 13125 31584
rect 12805 30496 13125 31520
rect 12805 30432 12813 30496
rect 12877 30432 12893 30496
rect 12957 30432 12973 30496
rect 13037 30432 13053 30496
rect 13117 30432 13125 30496
rect 12805 29408 13125 30432
rect 12805 29344 12813 29408
rect 12877 29344 12893 29408
rect 12957 29344 12973 29408
rect 13037 29344 13053 29408
rect 13117 29344 13125 29408
rect 12805 28320 13125 29344
rect 12805 28256 12813 28320
rect 12877 28256 12893 28320
rect 12957 28256 12973 28320
rect 13037 28256 13053 28320
rect 13117 28256 13125 28320
rect 12805 27232 13125 28256
rect 12805 27168 12813 27232
rect 12877 27168 12893 27232
rect 12957 27168 12973 27232
rect 13037 27168 13053 27232
rect 13117 27168 13125 27232
rect 12805 26144 13125 27168
rect 12805 26080 12813 26144
rect 12877 26080 12893 26144
rect 12957 26080 12973 26144
rect 13037 26080 13053 26144
rect 13117 26080 13125 26144
rect 12805 25056 13125 26080
rect 12805 24992 12813 25056
rect 12877 24992 12893 25056
rect 12957 24992 12973 25056
rect 13037 24992 13053 25056
rect 13117 24992 13125 25056
rect 12805 23968 13125 24992
rect 12805 23904 12813 23968
rect 12877 23904 12893 23968
rect 12957 23904 12973 23968
rect 13037 23904 13053 23968
rect 13117 23904 13125 23968
rect 12805 22880 13125 23904
rect 12805 22816 12813 22880
rect 12877 22816 12893 22880
rect 12957 22816 12973 22880
rect 13037 22816 13053 22880
rect 13117 22816 13125 22880
rect 12805 21792 13125 22816
rect 12805 21728 12813 21792
rect 12877 21728 12893 21792
rect 12957 21728 12973 21792
rect 13037 21728 13053 21792
rect 13117 21728 13125 21792
rect 12805 20704 13125 21728
rect 12805 20640 12813 20704
rect 12877 20640 12893 20704
rect 12957 20640 12973 20704
rect 13037 20640 13053 20704
rect 13117 20640 13125 20704
rect 12805 19616 13125 20640
rect 12805 19552 12813 19616
rect 12877 19552 12893 19616
rect 12957 19552 12973 19616
rect 13037 19552 13053 19616
rect 13117 19552 13125 19616
rect 12805 18528 13125 19552
rect 12805 18464 12813 18528
rect 12877 18464 12893 18528
rect 12957 18464 12973 18528
rect 13037 18464 13053 18528
rect 13117 18464 13125 18528
rect 12805 17440 13125 18464
rect 12805 17376 12813 17440
rect 12877 17376 12893 17440
rect 12957 17376 12973 17440
rect 13037 17376 13053 17440
rect 13117 17376 13125 17440
rect 12805 16352 13125 17376
rect 12805 16288 12813 16352
rect 12877 16288 12893 16352
rect 12957 16288 12973 16352
rect 13037 16288 13053 16352
rect 13117 16288 13125 16352
rect 12805 15264 13125 16288
rect 12805 15200 12813 15264
rect 12877 15200 12893 15264
rect 12957 15200 12973 15264
rect 13037 15200 13053 15264
rect 13117 15200 13125 15264
rect 12805 14176 13125 15200
rect 12805 14112 12813 14176
rect 12877 14112 12893 14176
rect 12957 14112 12973 14176
rect 13037 14112 13053 14176
rect 13117 14112 13125 14176
rect 12805 13088 13125 14112
rect 12805 13024 12813 13088
rect 12877 13024 12893 13088
rect 12957 13024 12973 13088
rect 13037 13024 13053 13088
rect 13117 13024 13125 13088
rect 12805 12000 13125 13024
rect 12805 11936 12813 12000
rect 12877 11936 12893 12000
rect 12957 11936 12973 12000
rect 13037 11936 13053 12000
rect 13117 11936 13125 12000
rect 12805 10912 13125 11936
rect 12805 10848 12813 10912
rect 12877 10848 12893 10912
rect 12957 10848 12973 10912
rect 13037 10848 13053 10912
rect 13117 10848 13125 10912
rect 12805 9824 13125 10848
rect 12805 9760 12813 9824
rect 12877 9760 12893 9824
rect 12957 9760 12973 9824
rect 13037 9760 13053 9824
rect 13117 9760 13125 9824
rect 12805 8736 13125 9760
rect 12805 8672 12813 8736
rect 12877 8672 12893 8736
rect 12957 8672 12973 8736
rect 13037 8672 13053 8736
rect 13117 8672 13125 8736
rect 12805 7648 13125 8672
rect 12805 7584 12813 7648
rect 12877 7584 12893 7648
rect 12957 7584 12973 7648
rect 13037 7584 13053 7648
rect 13117 7584 13125 7648
rect 12805 6560 13125 7584
rect 12805 6496 12813 6560
rect 12877 6496 12893 6560
rect 12957 6496 12973 6560
rect 13037 6496 13053 6560
rect 13117 6496 13125 6560
rect 12805 5472 13125 6496
rect 12805 5408 12813 5472
rect 12877 5408 12893 5472
rect 12957 5408 12973 5472
rect 13037 5408 13053 5472
rect 13117 5408 13125 5472
rect 12805 4384 13125 5408
rect 12805 4320 12813 4384
rect 12877 4320 12893 4384
rect 12957 4320 12973 4384
rect 13037 4320 13053 4384
rect 13117 4320 13125 4384
rect 12805 3296 13125 4320
rect 12805 3232 12813 3296
rect 12877 3232 12893 3296
rect 12957 3232 12973 3296
rect 13037 3232 13053 3296
rect 13117 3232 13125 3296
rect 12805 2208 13125 3232
rect 12805 2144 12813 2208
rect 12877 2144 12893 2208
rect 12957 2144 12973 2208
rect 13037 2144 13053 2208
rect 13117 2144 13125 2208
rect 12805 2128 13125 2144
rect 15770 47360 16091 47376
rect 15770 47296 15778 47360
rect 15842 47296 15858 47360
rect 15922 47296 15938 47360
rect 16002 47296 16018 47360
rect 16082 47296 16091 47360
rect 15770 46272 16091 47296
rect 15770 46208 15778 46272
rect 15842 46208 15858 46272
rect 15922 46208 15938 46272
rect 16002 46208 16018 46272
rect 16082 46208 16091 46272
rect 15770 45184 16091 46208
rect 15770 45120 15778 45184
rect 15842 45120 15858 45184
rect 15922 45120 15938 45184
rect 16002 45120 16018 45184
rect 16082 45120 16091 45184
rect 15770 44096 16091 45120
rect 15770 44032 15778 44096
rect 15842 44032 15858 44096
rect 15922 44032 15938 44096
rect 16002 44032 16018 44096
rect 16082 44032 16091 44096
rect 15770 43008 16091 44032
rect 15770 42944 15778 43008
rect 15842 42944 15858 43008
rect 15922 42944 15938 43008
rect 16002 42944 16018 43008
rect 16082 42944 16091 43008
rect 15770 41920 16091 42944
rect 15770 41856 15778 41920
rect 15842 41856 15858 41920
rect 15922 41856 15938 41920
rect 16002 41856 16018 41920
rect 16082 41856 16091 41920
rect 15770 40832 16091 41856
rect 15770 40768 15778 40832
rect 15842 40768 15858 40832
rect 15922 40768 15938 40832
rect 16002 40768 16018 40832
rect 16082 40768 16091 40832
rect 15770 39744 16091 40768
rect 15770 39680 15778 39744
rect 15842 39680 15858 39744
rect 15922 39680 15938 39744
rect 16002 39680 16018 39744
rect 16082 39680 16091 39744
rect 15770 38656 16091 39680
rect 15770 38592 15778 38656
rect 15842 38592 15858 38656
rect 15922 38592 15938 38656
rect 16002 38592 16018 38656
rect 16082 38592 16091 38656
rect 15770 37568 16091 38592
rect 15770 37504 15778 37568
rect 15842 37504 15858 37568
rect 15922 37504 15938 37568
rect 16002 37504 16018 37568
rect 16082 37504 16091 37568
rect 15770 36480 16091 37504
rect 15770 36416 15778 36480
rect 15842 36416 15858 36480
rect 15922 36416 15938 36480
rect 16002 36416 16018 36480
rect 16082 36416 16091 36480
rect 15770 35392 16091 36416
rect 15770 35328 15778 35392
rect 15842 35328 15858 35392
rect 15922 35328 15938 35392
rect 16002 35328 16018 35392
rect 16082 35328 16091 35392
rect 15770 34304 16091 35328
rect 15770 34240 15778 34304
rect 15842 34240 15858 34304
rect 15922 34240 15938 34304
rect 16002 34240 16018 34304
rect 16082 34240 16091 34304
rect 15770 33216 16091 34240
rect 15770 33152 15778 33216
rect 15842 33152 15858 33216
rect 15922 33152 15938 33216
rect 16002 33152 16018 33216
rect 16082 33152 16091 33216
rect 15770 32128 16091 33152
rect 15770 32064 15778 32128
rect 15842 32064 15858 32128
rect 15922 32064 15938 32128
rect 16002 32064 16018 32128
rect 16082 32064 16091 32128
rect 15770 31040 16091 32064
rect 15770 30976 15778 31040
rect 15842 30976 15858 31040
rect 15922 30976 15938 31040
rect 16002 30976 16018 31040
rect 16082 30976 16091 31040
rect 15770 29952 16091 30976
rect 15770 29888 15778 29952
rect 15842 29888 15858 29952
rect 15922 29888 15938 29952
rect 16002 29888 16018 29952
rect 16082 29888 16091 29952
rect 15770 28864 16091 29888
rect 15770 28800 15778 28864
rect 15842 28800 15858 28864
rect 15922 28800 15938 28864
rect 16002 28800 16018 28864
rect 16082 28800 16091 28864
rect 15770 27776 16091 28800
rect 15770 27712 15778 27776
rect 15842 27712 15858 27776
rect 15922 27712 15938 27776
rect 16002 27712 16018 27776
rect 16082 27712 16091 27776
rect 15770 26688 16091 27712
rect 15770 26624 15778 26688
rect 15842 26624 15858 26688
rect 15922 26624 15938 26688
rect 16002 26624 16018 26688
rect 16082 26624 16091 26688
rect 15770 25600 16091 26624
rect 15770 25536 15778 25600
rect 15842 25536 15858 25600
rect 15922 25536 15938 25600
rect 16002 25536 16018 25600
rect 16082 25536 16091 25600
rect 15770 24512 16091 25536
rect 15770 24448 15778 24512
rect 15842 24448 15858 24512
rect 15922 24448 15938 24512
rect 16002 24448 16018 24512
rect 16082 24448 16091 24512
rect 15770 23424 16091 24448
rect 15770 23360 15778 23424
rect 15842 23360 15858 23424
rect 15922 23360 15938 23424
rect 16002 23360 16018 23424
rect 16082 23360 16091 23424
rect 15770 22336 16091 23360
rect 15770 22272 15778 22336
rect 15842 22272 15858 22336
rect 15922 22272 15938 22336
rect 16002 22272 16018 22336
rect 16082 22272 16091 22336
rect 15770 21248 16091 22272
rect 15770 21184 15778 21248
rect 15842 21184 15858 21248
rect 15922 21184 15938 21248
rect 16002 21184 16018 21248
rect 16082 21184 16091 21248
rect 15770 20160 16091 21184
rect 15770 20096 15778 20160
rect 15842 20096 15858 20160
rect 15922 20096 15938 20160
rect 16002 20096 16018 20160
rect 16082 20096 16091 20160
rect 15770 19072 16091 20096
rect 15770 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15938 19072
rect 16002 19008 16018 19072
rect 16082 19008 16091 19072
rect 15770 17984 16091 19008
rect 15770 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15938 17984
rect 16002 17920 16018 17984
rect 16082 17920 16091 17984
rect 15770 16896 16091 17920
rect 15770 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15938 16896
rect 16002 16832 16018 16896
rect 16082 16832 16091 16896
rect 15770 15808 16091 16832
rect 15770 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15938 15808
rect 16002 15744 16018 15808
rect 16082 15744 16091 15808
rect 15770 14720 16091 15744
rect 15770 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15938 14720
rect 16002 14656 16018 14720
rect 16082 14656 16091 14720
rect 15770 13632 16091 14656
rect 15770 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15938 13632
rect 16002 13568 16018 13632
rect 16082 13568 16091 13632
rect 15770 12544 16091 13568
rect 15770 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15938 12544
rect 16002 12480 16018 12544
rect 16082 12480 16091 12544
rect 15770 11456 16091 12480
rect 15770 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15938 11456
rect 16002 11392 16018 11456
rect 16082 11392 16091 11456
rect 15770 10368 16091 11392
rect 15770 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15938 10368
rect 16002 10304 16018 10368
rect 16082 10304 16091 10368
rect 15770 9280 16091 10304
rect 15770 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15938 9280
rect 16002 9216 16018 9280
rect 16082 9216 16091 9280
rect 15770 8192 16091 9216
rect 15770 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15938 8192
rect 16002 8128 16018 8192
rect 16082 8128 16091 8192
rect 15770 7104 16091 8128
rect 15770 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15938 7104
rect 16002 7040 16018 7104
rect 16082 7040 16091 7104
rect 15770 6016 16091 7040
rect 15770 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15938 6016
rect 16002 5952 16018 6016
rect 16082 5952 16091 6016
rect 15770 4928 16091 5952
rect 15770 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15938 4928
rect 16002 4864 16018 4928
rect 16082 4864 16091 4928
rect 15770 3840 16091 4864
rect 15770 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15938 3840
rect 16002 3776 16018 3840
rect 16082 3776 16091 3840
rect 15770 2752 16091 3776
rect 15770 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15938 2752
rect 16002 2688 16018 2752
rect 16082 2688 16091 2752
rect 15770 2128 16091 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1644511149
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_175
timestamp 1644511149
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1644511149
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1644511149
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1644511149
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1644511149
transform 1 0 11316 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1644511149
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_66
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_83
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 1644511149
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_131
timestamp 1644511149
transform 1 0 13156 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1644511149
transform 1 0 15180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1644511149
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_63
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_72
timestamp 1644511149
transform 1 0 7728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1644511149
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1644511149
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_108
timestamp 1644511149
transform 1 0 11040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1644511149
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1644511149
transform 1 0 14352 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_151
timestamp 1644511149
transform 1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_158
timestamp 1644511149
transform 1 0 15640 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_170
timestamp 1644511149
transform 1 0 16744 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_182
timestamp 1644511149
transform 1 0 17848 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_35
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_41
timestamp 1644511149
transform 1 0 4876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1644511149
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1644511149
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_75
timestamp 1644511149
transform 1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_84
timestamp 1644511149
transform 1 0 8832 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1644511149
transform 1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1644511149
transform 1 0 10028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1644511149
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_116
timestamp 1644511149
transform 1 0 11776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp 1644511149
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_156
timestamp 1644511149
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1644511149
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1644511149
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1644511149
transform 1 0 6164 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp 1644511149
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_67
timestamp 1644511149
transform 1 0 7268 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_75
timestamp 1644511149
transform 1 0 8004 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1644511149
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_107
timestamp 1644511149
transform 1 0 10948 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_116
timestamp 1644511149
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_126
timestamp 1644511149
transform 1 0 12696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1644511149
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1644511149
transform 1 0 14720 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1644511149
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_166
timestamp 1644511149
transform 1 0 16376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_173
timestamp 1644511149
transform 1 0 17020 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_181
timestamp 1644511149
transform 1 0 17756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1644511149
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1644511149
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1644511149
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp 1644511149
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1644511149
transform 1 0 7912 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1644511149
transform 1 0 9016 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1644511149
transform 1 0 10120 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1644511149
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1644511149
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1644511149
transform 1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1644511149
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1644511149
transform 1 0 15456 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1644511149
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_173
timestamp 1644511149
transform 1 0 17020 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_179
timestamp 1644511149
transform 1 0 17572 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_187
timestamp 1644511149
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1644511149
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_100
timestamp 1644511149
transform 1 0 10304 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_112
timestamp 1644511149
transform 1 0 11408 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_116
timestamp 1644511149
transform 1 0 11776 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_151
timestamp 1644511149
transform 1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_175
timestamp 1644511149
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_187
timestamp 1644511149
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp 1644511149
transform 1 0 8004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1644511149
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1644511149
transform 1 0 11960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_122
timestamp 1644511149
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_126
timestamp 1644511149
transform 1 0 12696 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_138
timestamp 1644511149
transform 1 0 13800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1644511149
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1644511149
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1644511149
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_113
timestamp 1644511149
transform 1 0 11500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_117
timestamp 1644511149
transform 1 0 11868 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1644511149
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_132
timestamp 1644511149
transform 1 0 13248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1644511149
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1644511149
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_152
timestamp 1644511149
transform 1 0 15088 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_164
timestamp 1644511149
transform 1 0 16192 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_176
timestamp 1644511149
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1644511149
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 1644511149
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1644511149
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_76
timestamp 1644511149
transform 1 0 8096 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_88
timestamp 1644511149
transform 1 0 9200 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_100
timestamp 1644511149
transform 1 0 10304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1644511149
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_120
timestamp 1644511149
transform 1 0 12144 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_132
timestamp 1644511149
transform 1 0 13248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_140
timestamp 1644511149
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_146
timestamp 1644511149
transform 1 0 14536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 1644511149
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1644511149
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_6
timestamp 1644511149
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_18
timestamp 1644511149
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1644511149
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_43
timestamp 1644511149
transform 1 0 5060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1644511149
transform 1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1644511149
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_71
timestamp 1644511149
transform 1 0 7636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_102
timestamp 1644511149
transform 1 0 10488 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_108
timestamp 1644511149
transform 1 0 11040 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_116
timestamp 1644511149
transform 1 0 11776 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_128
timestamp 1644511149
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1644511149
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1644511149
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1644511149
transform 1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_73
timestamp 1644511149
transform 1 0 7820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_85
timestamp 1644511149
transform 1 0 8924 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_91
timestamp 1644511149
transform 1 0 9476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1644511149
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1644511149
transform 1 0 5428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1644511149
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_66
timestamp 1644511149
transform 1 0 7176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_118
timestamp 1644511149
transform 1 0 11960 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1644511149
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1644511149
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_33
timestamp 1644511149
transform 1 0 4140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_40
timestamp 1644511149
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_64
timestamp 1644511149
transform 1 0 6992 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_74
timestamp 1644511149
transform 1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1644511149
transform 1 0 9752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1644511149
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_134
timestamp 1644511149
transform 1 0 13432 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_141
timestamp 1644511149
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_148
timestamp 1644511149
transform 1 0 14720 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1644511149
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1644511149
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_47
timestamp 1644511149
transform 1 0 5428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1644511149
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1644511149
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1644511149
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_103
timestamp 1644511149
transform 1 0 10580 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_116
timestamp 1644511149
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_147
timestamp 1644511149
transform 1 0 14628 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_170
timestamp 1644511149
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_182
timestamp 1644511149
transform 1 0 17848 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_44
timestamp 1644511149
transform 1 0 5152 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_71
timestamp 1644511149
transform 1 0 7636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_79
timestamp 1644511149
transform 1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1644511149
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_100
timestamp 1644511149
transform 1 0 10304 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1644511149
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1644511149
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1644511149
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_61
timestamp 1644511149
transform 1 0 6716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1644511149
transform 1 0 9660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_101
timestamp 1644511149
transform 1 0 10396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_123
timestamp 1644511149
transform 1 0 12420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1644511149
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_149
timestamp 1644511149
transform 1 0 14812 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_171
timestamp 1644511149
transform 1 0 16836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1644511149
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_77
timestamp 1644511149
transform 1 0 8188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_84
timestamp 1644511149
transform 1 0 8832 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_94
timestamp 1644511149
transform 1 0 9752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_101
timestamp 1644511149
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1644511149
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_150
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_158
timestamp 1644511149
transform 1 0 15640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1644511149
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1644511149
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_168
timestamp 1644511149
transform 1 0 16560 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1644511149
transform 1 0 17480 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_89
timestamp 1644511149
transform 1 0 9292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_96
timestamp 1644511149
transform 1 0 9936 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1644511149
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_133
timestamp 1644511149
transform 1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_141
timestamp 1644511149
transform 1 0 14076 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1644511149
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_34
timestamp 1644511149
transform 1 0 4232 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_46
timestamp 1644511149
transform 1 0 5336 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_58
timestamp 1644511149
transform 1 0 6440 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_70
timestamp 1644511149
transform 1 0 7544 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1644511149
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_91
timestamp 1644511149
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1644511149
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1644511149
transform 1 0 10856 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_118
timestamp 1644511149
transform 1 0 11960 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 1644511149
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1644511149
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_160
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_172
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_180
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_186
timestamp 1644511149
transform 1 0 18216 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_23
timestamp 1644511149
transform 1 0 3220 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_28
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_37
timestamp 1644511149
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 1644511149
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1644511149
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1644511149
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_73
timestamp 1644511149
transform 1 0 7820 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_88
timestamp 1644511149
transform 1 0 9200 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1644511149
transform 1 0 10396 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_121
timestamp 1644511149
transform 1 0 12236 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_133
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_145
timestamp 1644511149
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1644511149
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1644511149
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1644511149
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_183
timestamp 1644511149
transform 1 0 17940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_19
timestamp 1644511149
transform 1 0 2852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1644511149
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_46
timestamp 1644511149
transform 1 0 5336 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_50
timestamp 1644511149
transform 1 0 5704 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1644511149
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_68
timestamp 1644511149
transform 1 0 7360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1644511149
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_108
timestamp 1644511149
transform 1 0 11040 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_116
timestamp 1644511149
transform 1 0 11776 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1644511149
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1644511149
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_145
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_157
timestamp 1644511149
transform 1 0 15548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_169
timestamp 1644511149
transform 1 0 16652 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_181
timestamp 1644511149
transform 1 0 17756 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1644511149
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_34
timestamp 1644511149
transform 1 0 4232 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1644511149
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1644511149
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1644511149
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_88
timestamp 1644511149
transform 1 0 9200 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1644511149
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1644511149
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_134
timestamp 1644511149
transform 1 0 13432 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_146
timestamp 1644511149
transform 1 0 14536 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 1644511149
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1644511149
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1644511149
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_179
timestamp 1644511149
transform 1 0 17572 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_187
timestamp 1644511149
transform 1 0 18308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_19
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_48
timestamp 1644511149
transform 1 0 5520 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_60
timestamp 1644511149
transform 1 0 6624 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_105
timestamp 1644511149
transform 1 0 10764 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_126
timestamp 1644511149
transform 1 0 12696 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_145
timestamp 1644511149
transform 1 0 14444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_152
timestamp 1644511149
transform 1 0 15088 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1644511149
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_38
timestamp 1644511149
transform 1 0 4600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1644511149
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_73
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_86
timestamp 1644511149
transform 1 0 9016 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1644511149
transform 1 0 9568 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_99
timestamp 1644511149
transform 1 0 10212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_103
timestamp 1644511149
transform 1 0 10580 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_131
timestamp 1644511149
transform 1 0 13156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_140
timestamp 1644511149
transform 1 0 13984 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1644511149
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_160
timestamp 1644511149
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 1644511149
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_45
timestamp 1644511149
transform 1 0 5244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1644511149
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_71
timestamp 1644511149
transform 1 0 7636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1644511149
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_103
timestamp 1644511149
transform 1 0 10580 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_108
timestamp 1644511149
transform 1 0 11040 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_120
timestamp 1644511149
transform 1 0 12144 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_129
timestamp 1644511149
transform 1 0 12972 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1644511149
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_166
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_175
timestamp 1644511149
transform 1 0 17204 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_182
timestamp 1644511149
transform 1 0 17848 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_6
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_18
timestamp 1644511149
transform 1 0 2760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_30
timestamp 1644511149
transform 1 0 3864 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_62
timestamp 1644511149
transform 1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1644511149
transform 1 0 7544 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1644511149
transform 1 0 8648 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_126
timestamp 1644511149
transform 1 0 12696 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_134
timestamp 1644511149
transform 1 0 13432 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_151
timestamp 1644511149
transform 1 0 14996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1644511149
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_174
timestamp 1644511149
transform 1 0 17112 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_186
timestamp 1644511149
transform 1 0 18216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_47
timestamp 1644511149
transform 1 0 5428 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_51
timestamp 1644511149
transform 1 0 5796 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_63
timestamp 1644511149
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_75
timestamp 1644511149
transform 1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_124
timestamp 1644511149
transform 1 0 12512 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_130
timestamp 1644511149
transform 1 0 13064 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_160
timestamp 1644511149
transform 1 0 15824 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_180
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1644511149
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_89
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_131
timestamp 1644511149
transform 1 0 13156 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1644511149
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_184
timestamp 1644511149
transform 1 0 18032 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_73
timestamp 1644511149
transform 1 0 7820 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1644511149
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1644511149
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_101
timestamp 1644511149
transform 1 0 10396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_108
timestamp 1644511149
transform 1 0 11040 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_120
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1644511149
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_149
timestamp 1644511149
transform 1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_162
timestamp 1644511149
transform 1 0 16008 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_186
timestamp 1644511149
transform 1 0 18216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_31
timestamp 1644511149
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_43
timestamp 1644511149
transform 1 0 5060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1644511149
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_61
timestamp 1644511149
transform 1 0 6716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_74
timestamp 1644511149
transform 1 0 7912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1644511149
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_87
timestamp 1644511149
transform 1 0 9108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_100
timestamp 1644511149
transform 1 0 10304 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1644511149
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_131
timestamp 1644511149
transform 1 0 13156 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_143
timestamp 1644511149
transform 1 0 14260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_155
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1644511149
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_46
timestamp 1644511149
transform 1 0 5336 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_54
timestamp 1644511149
transform 1 0 6072 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_107
timestamp 1644511149
transform 1 0 10948 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_127
timestamp 1644511149
transform 1 0 12788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1644511149
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_181
timestamp 1644511149
transform 1 0 17756 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_185
timestamp 1644511149
transform 1 0 18124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_24
timestamp 1644511149
transform 1 0 3312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_28
timestamp 1644511149
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_37
timestamp 1644511149
transform 1 0 4508 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1644511149
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_73
timestamp 1644511149
transform 1 0 7820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1644511149
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1644511149
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_117
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_129
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1644511149
transform 1 0 13524 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1644511149
transform 1 0 14628 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1644511149
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_175
timestamp 1644511149
transform 1 0 17204 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_182
timestamp 1644511149
transform 1 0 17848 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_11
timestamp 1644511149
transform 1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_17
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_35
timestamp 1644511149
transform 1 0 4324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_46
timestamp 1644511149
transform 1 0 5336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_60
timestamp 1644511149
transform 1 0 6624 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_88
timestamp 1644511149
transform 1 0 9200 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_108
timestamp 1644511149
transform 1 0 11040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_115
timestamp 1644511149
transform 1 0 11684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_127
timestamp 1644511149
transform 1 0 12788 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_148
timestamp 1644511149
transform 1 0 14720 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_160
timestamp 1644511149
transform 1 0 15824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_166
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_175
timestamp 1644511149
transform 1 0 17204 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_184
timestamp 1644511149
transform 1 0 18032 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_19
timestamp 1644511149
transform 1 0 2852 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_24
timestamp 1644511149
transform 1 0 3312 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 1644511149
transform 1 0 4048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1644511149
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_73
timestamp 1644511149
transform 1 0 7820 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1644511149
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_103
timestamp 1644511149
transform 1 0 10580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_116
timestamp 1644511149
transform 1 0 11776 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_120
timestamp 1644511149
transform 1 0 12144 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_147
timestamp 1644511149
transform 1 0 14628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_185
timestamp 1644511149
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_37
timestamp 1644511149
transform 1 0 4508 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_43
timestamp 1644511149
transform 1 0 5060 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_50
timestamp 1644511149
transform 1 0 5704 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_58
timestamp 1644511149
transform 1 0 6440 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_62
timestamp 1644511149
transform 1 0 6808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_69
timestamp 1644511149
transform 1 0 7452 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_75
timestamp 1644511149
transform 1 0 8004 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1644511149
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_90
timestamp 1644511149
transform 1 0 9384 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_102
timestamp 1644511149
transform 1 0 10488 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_114
timestamp 1644511149
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_126
timestamp 1644511149
transform 1 0 12696 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1644511149
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_156
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_160
timestamp 1644511149
transform 1 0 15824 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_166
timestamp 1644511149
transform 1 0 16376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_186
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_19
timestamp 1644511149
transform 1 0 2852 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_26
timestamp 1644511149
transform 1 0 3496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_34
timestamp 1644511149
transform 1 0 4232 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_46
timestamp 1644511149
transform 1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1644511149
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_67
timestamp 1644511149
transform 1 0 7268 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1644511149
transform 1 0 7912 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1644511149
transform 1 0 9016 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1644511149
transform 1 0 10120 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1644511149
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_129
timestamp 1644511149
transform 1 0 12972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_133
timestamp 1644511149
transform 1 0 13340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_153
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_159
timestamp 1644511149
transform 1 0 15732 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_186
timestamp 1644511149
transform 1 0 18216 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_11
timestamp 1644511149
transform 1 0 2116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1644511149
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_33
timestamp 1644511149
transform 1 0 4140 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_46
timestamp 1644511149
transform 1 0 5336 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_58
timestamp 1644511149
transform 1 0 6440 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_70
timestamp 1644511149
transform 1 0 7544 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1644511149
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_103
timestamp 1644511149
transform 1 0 10580 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_124
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1644511149
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_169
timestamp 1644511149
transform 1 0 16652 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_173
timestamp 1644511149
transform 1 0 17020 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_181
timestamp 1644511149
transform 1 0 17756 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_129
timestamp 1644511149
transform 1 0 12972 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_144
timestamp 1644511149
transform 1 0 14352 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_176
timestamp 1644511149
transform 1 0 17296 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_186
timestamp 1644511149
transform 1 0 18216 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_37
timestamp 1644511149
transform 1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_49
timestamp 1644511149
transform 1 0 5612 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_58
timestamp 1644511149
transform 1 0 6440 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_70
timestamp 1644511149
transform 1 0 7544 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1644511149
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1644511149
transform 1 0 9476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_105
timestamp 1644511149
transform 1 0 10764 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_110
timestamp 1644511149
transform 1 0 11224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_119
timestamp 1644511149
transform 1 0 12052 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_128
timestamp 1644511149
transform 1 0 12880 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 1644511149
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_148
timestamp 1644511149
transform 1 0 14720 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_162
timestamp 1644511149
transform 1 0 16008 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_183
timestamp 1644511149
transform 1 0 17940 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_43
timestamp 1644511149
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_61
timestamp 1644511149
transform 1 0 6716 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_76
timestamp 1644511149
transform 1 0 8096 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_88
timestamp 1644511149
transform 1 0 9200 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_98
timestamp 1644511149
transform 1 0 10120 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_129
timestamp 1644511149
transform 1 0 12972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_153
timestamp 1644511149
transform 1 0 15180 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 1644511149
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_174
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_186
timestamp 1644511149
transform 1 0 18216 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_35
timestamp 1644511149
transform 1 0 4324 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_44
timestamp 1644511149
transform 1 0 5152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_64
timestamp 1644511149
transform 1 0 6992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_73
timestamp 1644511149
transform 1 0 7820 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1644511149
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_91
timestamp 1644511149
transform 1 0 9476 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_111
timestamp 1644511149
transform 1 0 11316 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_124
timestamp 1644511149
transform 1 0 12512 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_7
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_19
timestamp 1644511149
transform 1 0 2852 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_31
timestamp 1644511149
transform 1 0 3956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1644511149
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1644511149
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_65
timestamp 1644511149
transform 1 0 7084 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_83
timestamp 1644511149
transform 1 0 8740 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1644511149
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_116
timestamp 1644511149
transform 1 0 11776 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_126
timestamp 1644511149
transform 1 0 12696 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_138
timestamp 1644511149
transform 1 0 13800 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_150
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1644511149
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_174
timestamp 1644511149
transform 1 0 17112 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_186
timestamp 1644511149
transform 1 0 18216 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_47
timestamp 1644511149
transform 1 0 5428 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_61
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_79
timestamp 1644511149
transform 1 0 8372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_89
timestamp 1644511149
transform 1 0 9292 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_98
timestamp 1644511149
transform 1 0 10120 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_106
timestamp 1644511149
transform 1 0 10856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_110
timestamp 1644511149
transform 1 0 11224 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_127
timestamp 1644511149
transform 1 0 12788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_144
timestamp 1644511149
transform 1 0 14352 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_156
timestamp 1644511149
transform 1 0 15456 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_168
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_180
timestamp 1644511149
transform 1 0 17664 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_188
timestamp 1644511149
transform 1 0 18400 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_37
timestamp 1644511149
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1644511149
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_63
timestamp 1644511149
transform 1 0 6900 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_77
timestamp 1644511149
transform 1 0 8188 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_89
timestamp 1644511149
transform 1 0 9292 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_101
timestamp 1644511149
transform 1 0 10396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1644511149
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1644511149
transform 1 0 12788 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1644511149
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1644511149
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_172
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_184
timestamp 1644511149
transform 1 0 18032 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_46
timestamp 1644511149
transform 1 0 5336 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_57
timestamp 1644511149
transform 1 0 6348 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_70
timestamp 1644511149
transform 1 0 7544 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1644511149
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_101
timestamp 1644511149
transform 1 0 10396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_113
timestamp 1644511149
transform 1 0 11500 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_126
timestamp 1644511149
transform 1 0 12696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_135
timestamp 1644511149
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_148
timestamp 1644511149
transform 1 0 14720 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_156
timestamp 1644511149
transform 1 0 15456 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_175
timestamp 1644511149
transform 1 0 17204 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_187
timestamp 1644511149
transform 1 0 18308 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_11
timestamp 1644511149
transform 1 0 2116 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_20
timestamp 1644511149
transform 1 0 2944 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_29
timestamp 1644511149
transform 1 0 3772 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_37
timestamp 1644511149
transform 1 0 4508 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_46
timestamp 1644511149
transform 1 0 5336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1644511149
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_154
timestamp 1644511149
transform 1 0 15272 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_174
timestamp 1644511149
transform 1 0 17112 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_186
timestamp 1644511149
transform 1 0 18216 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1644511149
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_56
timestamp 1644511149
transform 1 0 6256 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_68
timestamp 1644511149
transform 1 0 7360 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1644511149
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_89
timestamp 1644511149
transform 1 0 9292 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_127
timestamp 1644511149
transform 1 0 12788 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_147
timestamp 1644511149
transform 1 0 14628 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_156
timestamp 1644511149
transform 1 0 15456 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_180
timestamp 1644511149
transform 1 0 17664 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_188
timestamp 1644511149
transform 1 0 18400 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_88
timestamp 1644511149
transform 1 0 9200 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_94
timestamp 1644511149
transform 1 0 9752 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_98
timestamp 1644511149
transform 1 0 10120 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_155
timestamp 1644511149
transform 1 0 15364 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1644511149
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_174
timestamp 1644511149
transform 1 0 17112 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_189
timestamp 1644511149
transform 1 0 18492 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1644511149
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_33
timestamp 1644511149
transform 1 0 4140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_45
timestamp 1644511149
transform 1 0 5244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_57
timestamp 1644511149
transform 1 0 6348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_74
timestamp 1644511149
transform 1 0 7912 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1644511149
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_88
timestamp 1644511149
transform 1 0 9200 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_92
timestamp 1644511149
transform 1 0 9568 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_98
timestamp 1644511149
transform 1 0 10120 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_106
timestamp 1644511149
transform 1 0 10856 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_118
timestamp 1644511149
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_130
timestamp 1644511149
transform 1 0 13064 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 1644511149
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_157
timestamp 1644511149
transform 1 0 15548 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_11
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_20
timestamp 1644511149
transform 1 0 2944 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_28
timestamp 1644511149
transform 1 0 3680 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_36
timestamp 1644511149
transform 1 0 4416 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_42
timestamp 1644511149
transform 1 0 4968 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_46
timestamp 1644511149
transform 1 0 5336 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1644511149
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_61
timestamp 1644511149
transform 1 0 6716 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_68
timestamp 1644511149
transform 1 0 7360 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_76
timestamp 1644511149
transform 1 0 8096 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_86
timestamp 1644511149
transform 1 0 9016 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_101
timestamp 1644511149
transform 1 0 10396 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_109
timestamp 1644511149
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_117
timestamp 1644511149
transform 1 0 11868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_129
timestamp 1644511149
transform 1 0 12972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_141
timestamp 1644511149
transform 1 0 14076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_147
timestamp 1644511149
transform 1 0 14628 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_159
timestamp 1644511149
transform 1 0 15732 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_172
timestamp 1644511149
transform 1 0 16928 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_184
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_36
timestamp 1644511149
transform 1 0 4416 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_43
timestamp 1644511149
transform 1 0 5060 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_56
timestamp 1644511149
transform 1 0 6256 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_68
timestamp 1644511149
transform 1 0 7360 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_89
timestamp 1644511149
transform 1 0 9292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_100
timestamp 1644511149
transform 1 0 10304 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_110
timestamp 1644511149
transform 1 0 11224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_114
timestamp 1644511149
transform 1 0 11592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_120
timestamp 1644511149
transform 1 0 12144 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_127
timestamp 1644511149
transform 1 0 12788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_43
timestamp 1644511149
transform 1 0 5060 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1644511149
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_63
timestamp 1644511149
transform 1 0 6900 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_71
timestamp 1644511149
transform 1 0 7636 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_77
timestamp 1644511149
transform 1 0 8188 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_87
timestamp 1644511149
transform 1 0 9108 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_95
timestamp 1644511149
transform 1 0 9844 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_100
timestamp 1644511149
transform 1 0 10304 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1644511149
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_122
timestamp 1644511149
transform 1 0 12328 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_132
timestamp 1644511149
transform 1 0 13248 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_140
timestamp 1644511149
transform 1 0 13984 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_152
timestamp 1644511149
transform 1 0 15088 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_189
timestamp 1644511149
transform 1 0 18492 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_35
timestamp 1644511149
transform 1 0 4324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_49
timestamp 1644511149
transform 1 0 5612 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_69
timestamp 1644511149
transform 1 0 7452 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1644511149
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_90
timestamp 1644511149
transform 1 0 9384 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_96
timestamp 1644511149
transform 1 0 9936 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_101
timestamp 1644511149
transform 1 0 10396 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_129
timestamp 1644511149
transform 1 0 12972 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp 1644511149
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_146
timestamp 1644511149
transform 1 0 14536 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_162
timestamp 1644511149
transform 1 0 16008 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_174
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_186
timestamp 1644511149
transform 1 0 18216 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_35
timestamp 1644511149
transform 1 0 4324 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1644511149
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_63
timestamp 1644511149
transform 1 0 6900 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_67
timestamp 1644511149
transform 1 0 7268 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_72
timestamp 1644511149
transform 1 0 7728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_80
timestamp 1644511149
transform 1 0 8464 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_88
timestamp 1644511149
transform 1 0 9200 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_100
timestamp 1644511149
transform 1 0 10304 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1644511149
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_122
timestamp 1644511149
transform 1 0 12328 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_132
timestamp 1644511149
transform 1 0 13248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_140
timestamp 1644511149
transform 1 0 13984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_152
timestamp 1644511149
transform 1 0 15088 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_189
timestamp 1644511149
transform 1 0 18492 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_49
timestamp 1644511149
transform 1 0 5612 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_55
timestamp 1644511149
transform 1 0 6164 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_62
timestamp 1644511149
transform 1 0 6808 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_70
timestamp 1644511149
transform 1 0 7544 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_75
timestamp 1644511149
transform 1 0 8004 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_117
timestamp 1644511149
transform 1 0 11868 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_134
timestamp 1644511149
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1644511149
transform 1 0 14352 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_156
timestamp 1644511149
transform 1 0 15456 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_163
timestamp 1644511149
transform 1 0 16100 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_175
timestamp 1644511149
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_187
timestamp 1644511149
transform 1 0 18308 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_99
timestamp 1644511149
transform 1 0 10212 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_104
timestamp 1644511149
transform 1 0 10672 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_119
timestamp 1644511149
transform 1 0 12052 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_127
timestamp 1644511149
transform 1 0 12788 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_147
timestamp 1644511149
transform 1 0 14628 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1644511149
transform 1 0 16928 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_184
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_73
timestamp 1644511149
transform 1 0 7820 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_78
timestamp 1644511149
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_150
timestamp 1644511149
transform 1 0 14904 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_154
timestamp 1644511149
transform 1 0 15272 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_171
timestamp 1644511149
transform 1 0 16836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_183
timestamp 1644511149
transform 1 0 17940 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_13
timestamp 1644511149
transform 1 0 2300 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_25
timestamp 1644511149
transform 1 0 3404 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_37
timestamp 1644511149
transform 1 0 4508 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_46
timestamp 1644511149
transform 1 0 5336 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_95
timestamp 1644511149
transform 1 0 9844 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_107
timestamp 1644511149
transform 1 0 10948 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_144
timestamp 1644511149
transform 1 0 14352 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_175
timestamp 1644511149
transform 1 0 17204 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_187
timestamp 1644511149
transform 1 0 18308 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_32
timestamp 1644511149
transform 1 0 4048 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_39
timestamp 1644511149
transform 1 0 4692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_51
timestamp 1644511149
transform 1 0 5796 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_63
timestamp 1644511149
transform 1 0 6900 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_71
timestamp 1644511149
transform 1 0 7636 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_79
timestamp 1644511149
transform 1 0 8372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_101
timestamp 1644511149
transform 1 0 10396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_108
timestamp 1644511149
transform 1 0 11040 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_120
timestamp 1644511149
transform 1 0 12144 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_132
timestamp 1644511149
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_147
timestamp 1644511149
transform 1 0 14628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_164
timestamp 1644511149
transform 1 0 16192 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_176
timestamp 1644511149
transform 1 0 17296 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_188
timestamp 1644511149
transform 1 0 18400 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_11
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_20
timestamp 1644511149
transform 1 0 2944 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_35
timestamp 1644511149
transform 1 0 4324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_45
timestamp 1644511149
transform 1 0 5244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_61
timestamp 1644511149
transform 1 0 6716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_103
timestamp 1644511149
transform 1 0 10580 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_160
timestamp 1644511149
transform 1 0 15824 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_189
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1644511149
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_37
timestamp 1644511149
transform 1 0 4508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1644511149
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_56
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_61
timestamp 1644511149
transform 1 0 6716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_95
timestamp 1644511149
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_103
timestamp 1644511149
transform 1 0 10580 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_117
timestamp 1644511149
transform 1 0 11868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_124
timestamp 1644511149
transform 1 0 12512 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_136
timestamp 1644511149
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_23
timestamp 1644511149
transform 1 0 3220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_29
timestamp 1644511149
transform 1 0 3772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_46
timestamp 1644511149
transform 1 0 5336 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1644511149
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_61
timestamp 1644511149
transform 1 0 6716 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_78
timestamp 1644511149
transform 1 0 8280 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_85
timestamp 1644511149
transform 1 0 8924 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_97
timestamp 1644511149
transform 1 0 10028 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_106
timestamp 1644511149
transform 1 0 10856 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_129
timestamp 1644511149
transform 1 0 12972 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_143
timestamp 1644511149
transform 1 0 14260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_155
timestamp 1644511149
transform 1 0 15364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_189
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1644511149
transform 1 0 4048 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_44
timestamp 1644511149
transform 1 0 5152 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_61
timestamp 1644511149
transform 1 0 6716 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_75
timestamp 1644511149
transform 1 0 8004 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_98
timestamp 1644511149
transform 1 0 10120 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_108
timestamp 1644511149
transform 1 0 11040 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_119
timestamp 1644511149
transform 1 0 12052 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_126
timestamp 1644511149
transform 1 0 12696 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_132
timestamp 1644511149
transform 1 0 13248 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_136
timestamp 1644511149
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_157
timestamp 1644511149
transform 1 0 15548 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_169
timestamp 1644511149
transform 1 0 16652 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_181
timestamp 1644511149
transform 1 0 17756 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_43
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_47
timestamp 1644511149
transform 1 0 5428 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_52
timestamp 1644511149
transform 1 0 5888 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_73
timestamp 1644511149
transform 1 0 7820 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_86
timestamp 1644511149
transform 1 0 9016 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_96
timestamp 1644511149
transform 1 0 9936 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_107
timestamp 1644511149
transform 1 0 10948 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_120
timestamp 1644511149
transform 1 0 12144 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_144
timestamp 1644511149
transform 1 0 14352 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_155
timestamp 1644511149
transform 1 0 15364 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_162
timestamp 1644511149
transform 1 0 16008 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_189
timestamp 1644511149
transform 1 0 18492 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_58
timestamp 1644511149
transform 1 0 6440 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_72
timestamp 1644511149
transform 1 0 7728 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_80
timestamp 1644511149
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_100
timestamp 1644511149
transform 1 0 10304 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_108
timestamp 1644511149
transform 1 0 11040 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_114
timestamp 1644511149
transform 1 0 11592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_119
timestamp 1644511149
transform 1 0 12052 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_128
timestamp 1644511149
transform 1 0 12880 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_132
timestamp 1644511149
transform 1 0 13248 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1644511149
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_151
timestamp 1644511149
transform 1 0 14996 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_160
timestamp 1644511149
transform 1 0 15824 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_169
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_181
timestamp 1644511149
transform 1 0 17756 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_47
timestamp 1644511149
transform 1 0 5428 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1644511149
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_63
timestamp 1644511149
transform 1 0 6900 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_78
timestamp 1644511149
transform 1 0 8280 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_90
timestamp 1644511149
transform 1 0 9384 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_98
timestamp 1644511149
transform 1 0 10120 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_107
timestamp 1644511149
transform 1 0 10948 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_117
timestamp 1644511149
transform 1 0 11868 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_121
timestamp 1644511149
transform 1 0 12236 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_141
timestamp 1644511149
transform 1 0 14076 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_147
timestamp 1644511149
transform 1 0 14628 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1644511149
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_174
timestamp 1644511149
transform 1 0 17112 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_186
timestamp 1644511149
transform 1 0 18216 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_59
timestamp 1644511149
transform 1 0 6532 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_73
timestamp 1644511149
transform 1 0 7820 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_79
timestamp 1644511149
transform 1 0 8372 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_89
timestamp 1644511149
transform 1 0 9292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_101
timestamp 1644511149
transform 1 0 10396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_113
timestamp 1644511149
transform 1 0 11500 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_125
timestamp 1644511149
transform 1 0 12604 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_129
timestamp 1644511149
transform 1 0 12972 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_137
timestamp 1644511149
transform 1 0 13708 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_158
timestamp 1644511149
transform 1 0 15640 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_178
timestamp 1644511149
transform 1 0 17480 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_75
timestamp 1644511149
transform 1 0 8004 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_83
timestamp 1644511149
transform 1 0 8740 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_95
timestamp 1644511149
transform 1 0 9844 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_107
timestamp 1644511149
transform 1 0 10948 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_150
timestamp 1644511149
transform 1 0 14904 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_157
timestamp 1644511149
transform 1 0 15548 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1644511149
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_186
timestamp 1644511149
transform 1 0 18216 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_75
timestamp 1644511149
transform 1 0 8004 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_88
timestamp 1644511149
transform 1 0 9200 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_96
timestamp 1644511149
transform 1 0 9936 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_102
timestamp 1644511149
transform 1 0 10488 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1644511149
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_189
timestamp 1644511149
transform 1 0 18492 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_89
timestamp 1644511149
transform 1 0 9292 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_96
timestamp 1644511149
transform 1 0 9936 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_104
timestamp 1644511149
transform 1 0 10672 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_63
timestamp 1644511149
transform 1 0 6900 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_73
timestamp 1644511149
transform 1 0 7820 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_79
timestamp 1644511149
transform 1 0 8372 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_87
timestamp 1644511149
transform 1 0 9108 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_96
timestamp 1644511149
transform 1 0 9936 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_106
timestamp 1644511149
transform 1 0 10856 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_124
timestamp 1644511149
transform 1 0 12512 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_136
timestamp 1644511149
transform 1 0 13616 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_148
timestamp 1644511149
transform 1 0 14720 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_160
timestamp 1644511149
transform 1 0 15824 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_189
timestamp 1644511149
transform 1 0 18492 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_59
timestamp 1644511149
transform 1 0 6532 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_79
timestamp 1644511149
transform 1 0 8372 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_101
timestamp 1644511149
transform 1 0 10396 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_114
timestamp 1644511149
transform 1 0 11592 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_125
timestamp 1644511149
transform 1 0 12604 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_135
timestamp 1644511149
transform 1 0 13524 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_13
timestamp 1644511149
transform 1 0 2300 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_25
timestamp 1644511149
transform 1 0 3404 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_37
timestamp 1644511149
transform 1 0 4508 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_52
timestamp 1644511149
transform 1 0 5888 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_73
timestamp 1644511149
transform 1 0 7820 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_83
timestamp 1644511149
transform 1 0 8740 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_91
timestamp 1644511149
transform 1 0 9476 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_108
timestamp 1644511149
transform 1 0 11040 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_129
timestamp 1644511149
transform 1 0 12972 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_141
timestamp 1644511149
transform 1 0 14076 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_153
timestamp 1644511149
transform 1 0 15180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_165
timestamp 1644511149
transform 1 0 16284 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_189
timestamp 1644511149
transform 1 0 18492 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_47
timestamp 1644511149
transform 1 0 5428 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_64
timestamp 1644511149
transform 1 0 6992 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_73
timestamp 1644511149
transform 1 0 7820 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_80
timestamp 1644511149
transform 1 0 8464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_101
timestamp 1644511149
transform 1 0 10396 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_115
timestamp 1644511149
transform 1 0 11684 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_122
timestamp 1644511149
transform 1 0 12328 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_134
timestamp 1644511149
transform 1 0 13432 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_65
timestamp 1644511149
transform 1 0 7084 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_72
timestamp 1644511149
transform 1 0 7728 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_91
timestamp 1644511149
transform 1 0 9476 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_99
timestamp 1644511149
transform 1 0 10212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_116
timestamp 1644511149
transform 1 0 11776 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_128
timestamp 1644511149
transform 1 0 12880 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_140
timestamp 1644511149
transform 1 0 13984 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_152
timestamp 1644511149
transform 1 0 15088 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1644511149
transform 1 0 16192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_189
timestamp 1644511149
transform 1 0 18492 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_88
timestamp 1644511149
transform 1 0 9200 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_100
timestamp 1644511149
transform 1 0 10304 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_112
timestamp 1644511149
transform 1 0 11408 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_124
timestamp 1644511149
transform 1 0 12512 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1644511149
transform 1 0 13616 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_189
timestamp 1644511149
transform 1 0 18492 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_15
timestamp 1644511149
transform 1 0 2484 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1644511149
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_69
timestamp 1644511149
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1644511149
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_116
timestamp 1644511149
transform 1 0 11776 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_128
timestamp 1644511149
transform 1 0 12880 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_169
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_181
timestamp 1644511149
transform 1 0 17756 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_186
timestamp 1644511149
transform 1 0 18216 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 18860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 18860 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 18860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 18860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 18860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 18860 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 18860 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 18860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 18860 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 18860 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 18860 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 18860 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0459_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12052 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1644511149
transform -1 0 11132 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1644511149
transform -1 0 9936 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0462_
timestamp 1644511149
transform -1 0 9292 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463_
timestamp 1644511149
transform -1 0 8924 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0464_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7912 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0465_
timestamp 1644511149
transform -1 0 8280 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0466_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6808 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1644511149
transform -1 0 8004 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0468_
timestamp 1644511149
transform -1 0 6716 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0469_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7452 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0470_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0471_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8280 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0472_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8096 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0473_
timestamp 1644511149
transform 1 0 8372 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0474_
timestamp 1644511149
transform 1 0 9200 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0475_
timestamp 1644511149
transform 1 0 10764 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0476_
timestamp 1644511149
transform 1 0 6900 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0477_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _0478_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 11684 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1644511149
transform -1 0 13432 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0480_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0481_
timestamp 1644511149
transform 1 0 12144 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0482_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1644511149
transform 1 0 10672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1644511149
transform -1 0 10396 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1644511149
transform 1 0 10580 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1644511149
transform -1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0487_
timestamp 1644511149
transform 1 0 8464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1644511149
transform -1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1644511149
transform -1 0 9108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0490_
timestamp 1644511149
transform -1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0491_
timestamp 1644511149
transform -1 0 10212 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1644511149
transform -1 0 9200 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1644511149
transform -1 0 8280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0494_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9200 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0495_
timestamp 1644511149
transform -1 0 8464 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0496_
timestamp 1644511149
transform 1 0 8188 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _0497_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9200 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0498_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0499_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0500_
timestamp 1644511149
transform -1 0 9752 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0501_
timestamp 1644511149
transform 1 0 9568 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0502_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0503_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 15824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1644511149
transform 1 0 5612 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1644511149
transform 1 0 5060 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1644511149
transform 1 0 5060 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1644511149
transform 1 0 4968 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0509_
timestamp 1644511149
transform 1 0 5520 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1644511149
transform -1 0 5336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0511_
timestamp 1644511149
transform 1 0 5704 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1644511149
transform 1 0 4784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1644511149
transform -1 0 5796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0514_
timestamp 1644511149
transform -1 0 5888 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0515_
timestamp 1644511149
transform -1 0 5888 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0516_
timestamp 1644511149
transform -1 0 5152 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0517_
timestamp 1644511149
transform 1 0 5704 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0518_
timestamp 1644511149
transform -1 0 6256 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0519_
timestamp 1644511149
transform 1 0 6624 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0520_
timestamp 1644511149
transform -1 0 6256 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_2  _0521_
timestamp 1644511149
transform 1 0 4692 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0522_
timestamp 1644511149
transform 1 0 12788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0523_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12512 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0524_
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0525_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14720 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0526_
timestamp 1644511149
transform 1 0 13156 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0527_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12696 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0528_
timestamp 1644511149
transform -1 0 14628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0529_
timestamp 1644511149
transform 1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0530_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12788 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0531_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12052 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0532_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0533_
timestamp 1644511149
transform 1 0 9016 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1644511149
transform 1 0 10488 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0535_
timestamp 1644511149
transform -1 0 11040 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0536_
timestamp 1644511149
transform -1 0 12052 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1644511149
transform -1 0 11224 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0538_
timestamp 1644511149
transform 1 0 12420 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0539_
timestamp 1644511149
transform 1 0 13248 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0540_
timestamp 1644511149
transform 1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0541_
timestamp 1644511149
transform -1 0 15088 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0542_
timestamp 1644511149
transform 1 0 13064 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1644511149
transform -1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0544_
timestamp 1644511149
transform 1 0 13156 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1644511149
transform 1 0 15732 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0546_
timestamp 1644511149
transform -1 0 14628 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0547_
timestamp 1644511149
transform -1 0 13616 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0548_
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1644511149
transform 1 0 15640 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0550_
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0551_
timestamp 1644511149
transform -1 0 16192 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0552_
timestamp 1644511149
transform -1 0 15364 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0553_
timestamp 1644511149
transform 1 0 14444 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0554_
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0555_
timestamp 1644511149
transform -1 0 15180 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0556_
timestamp 1644511149
transform -1 0 14536 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1644511149
transform -1 0 14352 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0558_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0559_
timestamp 1644511149
transform 1 0 12420 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1644511149
transform -1 0 12972 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0561_
timestamp 1644511149
transform 1 0 14996 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0562_
timestamp 1644511149
transform 1 0 14444 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1644511149
transform -1 0 15548 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0564_
timestamp 1644511149
transform -1 0 15824 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0565_
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0566_
timestamp 1644511149
transform -1 0 14260 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1644511149
transform -1 0 13616 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0568_
timestamp 1644511149
transform -1 0 16652 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0569_
timestamp 1644511149
transform 1 0 15732 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0570_
timestamp 1644511149
transform -1 0 17112 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1644511149
transform -1 0 16192 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0572_
timestamp 1644511149
transform -1 0 15824 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1644511149
transform -1 0 14352 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0574_
timestamp 1644511149
transform 1 0 15088 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0575_
timestamp 1644511149
transform 1 0 15640 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0577_
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1644511149
transform -1 0 15732 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0579_
timestamp 1644511149
transform -1 0 17756 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0580_
timestamp 1644511149
transform -1 0 16836 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0581_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0582_
timestamp 1644511149
transform -1 0 18216 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0583_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0584_
timestamp 1644511149
transform 1 0 15272 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0585_
timestamp 1644511149
transform 1 0 12052 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0586_
timestamp 1644511149
transform -1 0 17940 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0587_
timestamp 1644511149
transform 1 0 17296 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0588_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0589_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0590_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1644511149
transform 1 0 17480 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0592_
timestamp 1644511149
transform -1 0 17112 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0594_
timestamp 1644511149
transform 1 0 14996 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0595_
timestamp 1644511149
transform 1 0 15916 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0596_
timestamp 1644511149
transform -1 0 17204 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1644511149
transform -1 0 17204 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1644511149
transform -1 0 16376 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0599_
timestamp 1644511149
transform -1 0 18032 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1644511149
transform 1 0 17572 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0601_
timestamp 1644511149
transform 1 0 13156 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1644511149
transform -1 0 13616 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0603_
timestamp 1644511149
transform -1 0 16560 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0604_
timestamp 1644511149
transform -1 0 16376 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0605_
timestamp 1644511149
transform 1 0 14260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0606_
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0607_
timestamp 1644511149
transform -1 0 16100 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0608_
timestamp 1644511149
transform 1 0 14536 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0609_
timestamp 1644511149
transform 1 0 9568 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1644511149
transform -1 0 11776 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0611_
timestamp 1644511149
transform 1 0 15180 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0612_
timestamp 1644511149
transform -1 0 17112 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0613_
timestamp 1644511149
transform 1 0 15548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0614_
timestamp 1644511149
transform 1 0 15548 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1644511149
transform -1 0 16928 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0616_
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1644511149
transform 1 0 17572 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0618_
timestamp 1644511149
transform 1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0619_
timestamp 1644511149
transform 1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0620_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1644511149
transform 1 0 17204 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0622_
timestamp 1644511149
transform -1 0 16008 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0624_
timestamp 1644511149
transform -1 0 12788 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0625_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0626_
timestamp 1644511149
transform -1 0 12696 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0627_
timestamp 1644511149
transform -1 0 11960 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0628_
timestamp 1644511149
transform -1 0 12972 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1644511149
transform 1 0 12144 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0630_
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0631_
timestamp 1644511149
transform -1 0 11960 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0632_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1644511149
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1644511149
transform 1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0635_
timestamp 1644511149
transform -1 0 10856 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1644511149
transform 1 0 10212 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0637_
timestamp 1644511149
transform -1 0 10764 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0639_
timestamp 1644511149
transform -1 0 10856 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 1644511149
transform 1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0641_
timestamp 1644511149
transform 1 0 10856 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1644511149
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0643_
timestamp 1644511149
transform 1 0 11316 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1644511149
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1644511149
transform -1 0 12880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0646_
timestamp 1644511149
transform 1 0 13064 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0647_
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0648_
timestamp 1644511149
transform -1 0 13616 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0649_
timestamp 1644511149
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0650_
timestamp 1644511149
transform 1 0 12972 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0651_
timestamp 1644511149
transform -1 0 14996 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0652_
timestamp 1644511149
transform -1 0 15088 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0653_
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0654_
timestamp 1644511149
transform -1 0 14352 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0655_
timestamp 1644511149
transform 1 0 13524 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1644511149
transform 1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0657_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0658_
timestamp 1644511149
transform -1 0 5336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0659_
timestamp 1644511149
transform 1 0 6164 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0660_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 5888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0661_
timestamp 1644511149
transform -1 0 6716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0662_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0663_
timestamp 1644511149
transform 1 0 5152 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0664_
timestamp 1644511149
transform 1 0 5244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0665_
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0666_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0667_
timestamp 1644511149
transform 1 0 7360 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0668_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0669_
timestamp 1644511149
transform -1 0 8464 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0670_
timestamp 1644511149
transform -1 0 7452 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0671_
timestamp 1644511149
transform -1 0 10856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0672_
timestamp 1644511149
transform -1 0 8188 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0673_
timestamp 1644511149
transform -1 0 7544 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0674_
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0675_
timestamp 1644511149
transform -1 0 8188 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0676_
timestamp 1644511149
transform -1 0 5888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0677_
timestamp 1644511149
transform 1 0 6808 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0678_
timestamp 1644511149
transform -1 0 6900 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0679_
timestamp 1644511149
transform 1 0 7268 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0680_
timestamp 1644511149
transform -1 0 6808 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1644511149
transform -1 0 7268 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0682_
timestamp 1644511149
transform 1 0 5796 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0683_
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0684_
timestamp 1644511149
transform 1 0 11684 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0685_
timestamp 1644511149
transform -1 0 12788 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0686_
timestamp 1644511149
transform -1 0 17572 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1644511149
transform 1 0 16744 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0688_
timestamp 1644511149
transform 1 0 14260 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1644511149
transform 1 0 14720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1644511149
transform 1 0 15088 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1644511149
transform 1 0 15824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0692_
timestamp 1644511149
transform -1 0 14536 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 1644511149
transform -1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0694_
timestamp 1644511149
transform -1 0 16376 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0695_
timestamp 1644511149
transform 1 0 15364 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0696_
timestamp 1644511149
transform -1 0 13432 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1644511149
transform 1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0698_
timestamp 1644511149
transform 1 0 13156 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 1644511149
transform -1 0 14076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0700_
timestamp 1644511149
transform 1 0 13616 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1644511149
transform -1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0702_
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0703_
timestamp 1644511149
transform 1 0 10580 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0704_
timestamp 1644511149
transform -1 0 12052 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0705_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12696 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0706_
timestamp 1644511149
transform -1 0 13248 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0707_
timestamp 1644511149
transform 1 0 11684 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0708_
timestamp 1644511149
transform -1 0 10396 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0709_
timestamp 1644511149
transform -1 0 11132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0710_
timestamp 1644511149
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0711_
timestamp 1644511149
transform 1 0 7820 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0712_
timestamp 1644511149
transform 1 0 11684 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0713_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0714_
timestamp 1644511149
transform -1 0 9384 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0715_
timestamp 1644511149
transform -1 0 8464 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0716_
timestamp 1644511149
transform 1 0 8004 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0717_
timestamp 1644511149
transform 1 0 8832 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0718_
timestamp 1644511149
transform -1 0 10120 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0719_
timestamp 1644511149
transform 1 0 8280 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0720_
timestamp 1644511149
transform 1 0 10672 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_2  _0721_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0722_
timestamp 1644511149
transform 1 0 9844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0723_
timestamp 1644511149
transform 1 0 9660 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1644511149
transform 1 0 10488 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0725_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9384 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0726_
timestamp 1644511149
transform 1 0 10120 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0727_
timestamp 1644511149
transform 1 0 9384 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0728_
timestamp 1644511149
transform 1 0 9936 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0729_
timestamp 1644511149
transform -1 0 10304 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0730_
timestamp 1644511149
transform 1 0 10488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _0731_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 11224 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0732_
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0733_
timestamp 1644511149
transform 1 0 9108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0734_
timestamp 1644511149
transform -1 0 11868 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0735_
timestamp 1644511149
transform -1 0 10396 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0736_
timestamp 1644511149
transform 1 0 9476 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0737_
timestamp 1644511149
transform 1 0 10764 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0738_
timestamp 1644511149
transform -1 0 10856 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0739_
timestamp 1644511149
transform -1 0 10580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0740_
timestamp 1644511149
transform 1 0 9292 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0741_
timestamp 1644511149
transform 1 0 9660 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0742_
timestamp 1644511149
transform 1 0 10672 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0743_
timestamp 1644511149
transform -1 0 9936 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0744_
timestamp 1644511149
transform 1 0 10304 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0745_
timestamp 1644511149
transform -1 0 10488 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0746_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10856 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0747_
timestamp 1644511149
transform 1 0 12420 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0748_
timestamp 1644511149
transform 1 0 11684 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0749_
timestamp 1644511149
transform 1 0 11960 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0750_
timestamp 1644511149
transform 1 0 10672 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0751_
timestamp 1644511149
transform -1 0 10948 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0752_
timestamp 1644511149
transform 1 0 11408 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0753_
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0754_
timestamp 1644511149
transform -1 0 11868 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0755_
timestamp 1644511149
transform 1 0 11684 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0756_
timestamp 1644511149
transform -1 0 12604 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0757_
timestamp 1644511149
transform 1 0 11868 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0758_
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0759_
timestamp 1644511149
transform 1 0 12972 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0760_
timestamp 1644511149
transform 1 0 13892 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0761_
timestamp 1644511149
transform -1 0 14720 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0762_
timestamp 1644511149
transform -1 0 8096 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0763_
timestamp 1644511149
transform -1 0 15456 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 1644511149
transform -1 0 13340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0765_
timestamp 1644511149
transform -1 0 14628 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0766_
timestamp 1644511149
transform -1 0 14628 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0767_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0768_
timestamp 1644511149
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0769_
timestamp 1644511149
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0770_
timestamp 1644511149
transform -1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0771_
timestamp 1644511149
transform -1 0 6716 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0772_
timestamp 1644511149
transform 1 0 12880 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0773_
timestamp 1644511149
transform -1 0 7820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0774_
timestamp 1644511149
transform -1 0 7636 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0775_
timestamp 1644511149
transform -1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0776_
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0777_
timestamp 1644511149
transform 1 0 7176 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0778_
timestamp 1644511149
transform -1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0779_
timestamp 1644511149
transform 1 0 5888 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0780_
timestamp 1644511149
transform -1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_2  _0781_
timestamp 1644511149
transform 1 0 6532 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1644511149
transform -1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0783_
timestamp 1644511149
transform -1 0 8832 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0784_
timestamp 1644511149
transform -1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0785_
timestamp 1644511149
transform -1 0 7268 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0786_
timestamp 1644511149
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0787_
timestamp 1644511149
transform -1 0 8004 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0788_
timestamp 1644511149
transform 1 0 7544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0789_
timestamp 1644511149
transform -1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0790_
timestamp 1644511149
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _0791_
timestamp 1644511149
transform -1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0792_
timestamp 1644511149
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0793_
timestamp 1644511149
transform -1 0 8372 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0794_
timestamp 1644511149
transform -1 0 7176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0795_
timestamp 1644511149
transform -1 0 7820 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0796_
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0797_
timestamp 1644511149
transform 1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0798_
timestamp 1644511149
transform 1 0 6808 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0799_
timestamp 1644511149
transform -1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0800_
timestamp 1644511149
transform 1 0 6900 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0801_
timestamp 1644511149
transform -1 0 6440 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0802_
timestamp 1644511149
transform -1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0803_
timestamp 1644511149
transform -1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0804_
timestamp 1644511149
transform -1 0 5796 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0805_
timestamp 1644511149
transform 1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0806_
timestamp 1644511149
transform -1 0 4784 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0807_
timestamp 1644511149
transform 1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0808_
timestamp 1644511149
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0809_
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0810_
timestamp 1644511149
transform 1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0811_
timestamp 1644511149
transform -1 0 6440 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0812_
timestamp 1644511149
transform 1 0 5152 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0814_
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0815_
timestamp 1644511149
transform -1 0 5612 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0816_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 5152 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0817_
timestamp 1644511149
transform -1 0 5336 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1644511149
transform 1 0 4968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0819_
timestamp 1644511149
transform -1 0 5060 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0820_
timestamp 1644511149
transform -1 0 14720 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0821_
timestamp 1644511149
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0822_
timestamp 1644511149
transform -1 0 5888 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0823_
timestamp 1644511149
transform -1 0 12696 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1644511149
transform -1 0 12512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0825_
timestamp 1644511149
transform -1 0 13616 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0826_
timestamp 1644511149
transform -1 0 13156 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0827_
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0828_
timestamp 1644511149
transform 1 0 4140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0829_
timestamp 1644511149
transform -1 0 5244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0830_
timestamp 1644511149
transform -1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0831_
timestamp 1644511149
transform 1 0 4968 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0832_
timestamp 1644511149
transform 1 0 11408 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0833_
timestamp 1644511149
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0834_
timestamp 1644511149
transform -1 0 4508 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0835_
timestamp 1644511149
transform -1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0836_
timestamp 1644511149
transform 1 0 2576 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0837_
timestamp 1644511149
transform 1 0 3312 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0838_
timestamp 1644511149
transform -1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0839_
timestamp 1644511149
transform 1 0 3864 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0840_
timestamp 1644511149
transform -1 0 4048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_2  _0841_
timestamp 1644511149
transform 1 0 3404 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 1644511149
transform -1 0 3312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1644511149
transform -1 0 4324 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0844_
timestamp 1644511149
transform 1 0 2392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0845_
timestamp 1644511149
transform 1 0 2668 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 1644511149
transform 1 0 3680 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0847_
timestamp 1644511149
transform 1 0 3772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0848_
timestamp 1644511149
transform -1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0849_
timestamp 1644511149
transform 1 0 2392 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0850_
timestamp 1644511149
transform 1 0 2944 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0851_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4508 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0852_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3496 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0853_
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0854_
timestamp 1644511149
transform -1 0 4140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0855_
timestamp 1644511149
transform 1 0 2668 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0856_
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 1644511149
transform -1 0 3312 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0858_
timestamp 1644511149
transform 1 0 3312 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0859_
timestamp 1644511149
transform 1 0 4140 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0860_
timestamp 1644511149
transform 1 0 3772 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0861_
timestamp 1644511149
transform 1 0 2300 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0862_
timestamp 1644511149
transform -1 0 3680 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0863_
timestamp 1644511149
transform -1 0 4140 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0864_
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1644511149
transform 1 0 4784 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0866_
timestamp 1644511149
transform -1 0 4324 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0867_
timestamp 1644511149
transform -1 0 4048 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0868_
timestamp 1644511149
transform -1 0 3312 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0869_
timestamp 1644511149
transform 1 0 2208 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0870_
timestamp 1644511149
transform -1 0 4416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0871_
timestamp 1644511149
transform 1 0 2668 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0872_
timestamp 1644511149
transform 1 0 2300 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0873_
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0874_
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0875_
timestamp 1644511149
transform 1 0 2852 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0876_
timestamp 1644511149
transform 1 0 3680 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0877_
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 1644511149
transform 1 0 4416 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0879_
timestamp 1644511149
transform -1 0 5244 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0880_
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1644511149
transform -1 0 5888 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0882_
timestamp 1644511149
transform 1 0 5520 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0883_
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0884_
timestamp 1644511149
transform -1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0885_
timestamp 1644511149
transform -1 0 7084 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0886_
timestamp 1644511149
transform -1 0 6716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0887_
timestamp 1644511149
transform -1 0 7820 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0888_
timestamp 1644511149
transform -1 0 6532 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0889_
timestamp 1644511149
transform -1 0 5888 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1644511149
transform 1 0 6992 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0891_
timestamp 1644511149
transform -1 0 7084 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0892_
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0893_
timestamp 1644511149
transform -1 0 8372 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1644511149
transform -1 0 8464 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0895_
timestamp 1644511149
transform 1 0 8188 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0896_
timestamp 1644511149
transform 1 0 8096 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0897_
timestamp 1644511149
transform -1 0 9292 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0898_
timestamp 1644511149
transform -1 0 9200 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0899_
timestamp 1644511149
transform -1 0 10212 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0900_
timestamp 1644511149
transform 1 0 8924 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0901_
timestamp 1644511149
transform -1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0902_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7636 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0903_
timestamp 1644511149
transform 1 0 7544 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0904_
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0905_
timestamp 1644511149
transform -1 0 9384 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0906_
timestamp 1644511149
transform -1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1644511149
transform 1 0 10028 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0908_
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0909_
timestamp 1644511149
transform 1 0 11408 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0910_
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0911_
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1644511149
transform 1 0 10764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0913_
timestamp 1644511149
transform 1 0 10580 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1644511149
transform -1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0915_
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0916_
timestamp 1644511149
transform -1 0 10396 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0917_
timestamp 1644511149
transform 1 0 11408 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0918_
timestamp 1644511149
transform -1 0 11040 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0919_
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0920_
timestamp 1644511149
transform 1 0 8648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _0921_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1644511149
transform 1 0 9844 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1644511149
transform 1 0 11316 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1644511149
transform -1 0 12972 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1644511149
transform -1 0 14628 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1644511149
transform -1 0 15548 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1644511149
transform 1 0 13892 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1644511149
transform -1 0 15272 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1644511149
transform -1 0 14628 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1644511149
transform -1 0 15640 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1644511149
transform 1 0 12880 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1644511149
transform 1 0 14720 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1644511149
transform 1 0 16008 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1644511149
transform 1 0 14720 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1644511149
transform 1 0 15364 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1644511149
transform 1 0 14720 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1644511149
transform -1 0 17388 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1644511149
transform 1 0 16192 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1644511149
transform 1 0 16744 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1644511149
transform 1 0 16744 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1644511149
transform -1 0 14996 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1644511149
transform 1 0 11316 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1644511149
transform -1 0 15824 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1644511149
transform -1 0 17664 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1644511149
transform -1 0 17480 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1644511149
transform 1 0 15364 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1644511149
transform -1 0 16744 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1644511149
transform 1 0 14720 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1644511149
transform 1 0 10948 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1644511149
transform 1 0 9568 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1644511149
transform 1 0 9476 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1644511149
transform 1 0 9568 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1644511149
transform 1 0 11408 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1644511149
transform -1 0 13156 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1644511149
transform -1 0 13616 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1644511149
transform 1 0 11868 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1644511149
transform 1 0 11592 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1644511149
transform -1 0 7820 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1644511149
transform 1 0 4416 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1644511149
transform -1 0 6992 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1644511149
transform -1 0 8740 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1644511149
transform 1 0 6900 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1644511149
transform 1 0 6440 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1644511149
transform 1 0 4416 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1644511149
transform -1 0 12972 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1644511149
transform -1 0 17204 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1644511149
transform 1 0 13984 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1644511149
transform -1 0 15456 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1644511149
transform 1 0 13984 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1644511149
transform -1 0 15180 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1644511149
transform 1 0 12052 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1644511149
transform -1 0 14904 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1644511149
transform -1 0 15548 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1644511149
transform -1 0 8556 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0986_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9108 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1644511149
transform 1 0 9108 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1644511149
transform -1 0 11040 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1644511149
transform -1 0 12972 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1644511149
transform -1 0 15180 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1644511149
transform -1 0 13432 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1644511149
transform 1 0 6992 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0997_
timestamp 1644511149
transform 1 0 8096 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1644511149
transform 1 0 6992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1644511149
transform 1 0 3956 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1644511149
transform 1 0 11224 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1644511149
transform 1 0 12236 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1644511149
transform 1 0 3864 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1644511149
transform 1 0 3864 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1644511149
transform 1 0 3864 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1644511149
transform 1 0 3864 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1644511149
transform -1 0 13432 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1644511149
transform 1 0 5244 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1644511149
transform 1 0 4968 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1644511149
transform 1 0 5520 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1644511149
transform -1 0 7820 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1644511149
transform 1 0 6900 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1644511149
transform 1 0 6992 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1644511149
transform 1 0 8188 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1644511149
transform 1 0 8372 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1644511149
transform 1 0 9568 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1644511149
transform -1 0 10948 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1644511149
transform 1 0 9292 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1644511149
transform -1 0 11040 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1644511149
transform 1 0 9108 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1029__12 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1030__13
timestamp 1644511149
transform -1 0 11776 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1031__14
timestamp 1644511149
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1032__15
timestamp 1644511149
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1644511149
transform 1 0 17848 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12512 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1644511149
transform 1 0 11868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform -1 0 10672 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clk
timestamp 1644511149
transform -1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clk
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clk
timestamp 1644511149
transform -1 0 8280 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clk
timestamp 1644511149
transform 1 0 12420 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clk
timestamp 1644511149
transform -1 0 9752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clk
timestamp 1644511149
transform -1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clk
timestamp 1644511149
transform 1 0 14444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clk
timestamp 1644511149
transform -1 0 14444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clk
timestamp 1644511149
transform -1 0 7728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clk
timestamp 1644511149
transform -1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clk
timestamp 1644511149
transform 1 0 13616 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clk
timestamp 1644511149
transform -1 0 13708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 17940 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 17940 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1644511149
transform 1 0 1748 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1644511149
transform 1 0 17848 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1644511149
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1644511149
transform -1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1644511149
transform -1 0 16192 0 -1 23936
box -38 -48 406 592
<< labels >>
rlabel metal3 s 19200 31968 20000 32088 6 clk
port 0 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 enc0_a
port 1 nsew signal input
rlabel metal3 s 19200 40808 20000 40928 6 enc0_b
port 2 nsew signal input
rlabel metal3 s 19200 14288 20000 14408 6 enc1_a
port 3 nsew signal input
rlabel metal2 s 2594 49200 2650 50000 6 enc1_b
port 4 nsew signal input
rlabel metal2 s 18 0 74 800 6 enc2_a
port 5 nsew signal input
rlabel metal3 s 19200 5448 20000 5568 6 enc2_b
port 6 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_oeb[0]
port 7 nsew signal tristate
rlabel metal2 s 10966 49200 11022 50000 6 io_oeb[1]
port 8 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 io_oeb[2]
port 9 nsew signal tristate
rlabel metal3 s 0 17688 800 17808 6 io_oeb[3]
port 10 nsew signal tristate
rlabel metal2 s 19338 49200 19394 50000 6 pwm0_out
port 11 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 pwm1_out
port 12 nsew signal tristate
rlabel metal3 s 0 26528 800 26648 6 pwm2_out
port 13 nsew signal tristate
rlabel metal3 s 0 44208 800 44328 6 reset
port 14 nsew signal input
rlabel metal3 s 19200 23128 20000 23248 6 sync
port 15 nsew signal tristate
rlabel metal4 s 3910 2128 4230 47376 6 vccd1
port 16 nsew power input
rlabel metal4 s 9840 2128 10160 47376 6 vccd1
port 16 nsew power input
rlabel metal4 s 15771 2128 16091 47376 6 vccd1
port 16 nsew power input
rlabel metal4 s 6874 2128 7194 47376 6 vssd1
port 17 nsew ground input
rlabel metal4 s 12805 2128 13125 47376 6 vssd1
port 17 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 20000 50000
<< end >>
